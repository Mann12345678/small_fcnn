library ieee;
use ieee.std_logic_1164.all;

entity layer_1 is
port ( 
       clk : in std_logic;
       Layer1_input : in std_logic_vector(4095 downto 0); ------------16 neuron
       Layer1_output : out std_logic_vector(255 downto 0)
       );
end entity;
    
architecture structure of layer_1 is 

component Neu_Ron is 
generic( N : integer := 4);
port ( clk : in std_logic; 
       inputs : in std_logic_vector( ((N*16)-1) downto 0);
       weights : in std_logic_vector( ((N*16)-1) downto 0);
       Bias : in std_logic_vector(15 downto 0);
       weighted_sum : out std_logic_vector(15 downto 0);
       neuron_output :out  std_logic_vector(15 downto 0)
      );
end component;

type weight_array is array (0 to 15) of std_logic_vector(4095 downto 0);
signal weight : weight_array := (
("0010100101000101001100001101101110101000111000100010110110000001101100010110011100100110001101100010101101001101101010000110010110101000010010001010010101001010101100001011001000100110000101010011001110110111101001101001100110100111000011000010011110010111101100100011101110100100011001110001100110000000101100010110110010110010001001110010100011110110001011000000111010010001010001110010110010011001101100001011001110100111111011010010111000011101001011001001000110110001011010101010110100001111001011101110110110110000001001100010010101110011101011000110100110110000000100000010001011100111101011110100001110011110111011110010111011010000101100001110000010011011000000001010101001100011001010001001011100110001011110011010100100000011001001110110001010101101111010101011000000001010001011101101110000011000011101101010101010011010101100010001000110101101110100110010110101010101001100000110000110101000110101111010101111010101101011010111101110101100010110100011000000010001001011110110010110101001000101010010100110101110101011001111110000101111010100011010110111110000101011011001110000110000000101010011000001011111001011011001100000110000101100010010110110000000101011010000010100101110010110011010100000001011001100010101011000101110010000011001101010000000101011100101110110110000010000000011000100001110101100001101111110101111011001001010101101001000101011010001111100110000111011010011000011000011001010111100110000100111111110100010110010000100001100001111010000011010010100101010111000001110001011011001000010101011011111010010101100101111001100000110011010100111001110101011000101101001001100001011011000101101110011100010010010011010101010001110000110101100111011100010110100100010101011011110110000101000101101110010111101100101100111111000010110101110101010000010010101110010100000110101100000110000100001011010010011110010101010101000000100110000001011111011000000110101101011111010110110100000011111101010011100101101101011100101001110101110010011110011000111111110001011101000110010101011000100010010111111010110101011101000101100101100011100011010110001010001001011001100111110101101101000100010010100010101000111000000110010101110010000001010101001011101101010011000101000101100110100110011000010101101101001101001001010110000011010101010110101011111001001111101100100110000010000000011000000010101001011001000011000011110101110010011000011100100101011001101111110101100011101111001101011000011001100101000011110110001000010110010100100101001101011100000000010101111111101110010110110101101101011000001000100101111000111110010111001011110001010010001000000101001111011101010111010100110001011110011110100101110110001111011000100000010001010101111011000100001011011110010110010001111101010011011110110101100110010110010011110011001101001010001101100011111110000111010101101000011001011101110111100010111110011001010100110011111001011011111010110110000101010001010110001110011001011111000100010110010101000111010111000000110101011110011011000101001011011111010010000101111101011111010010010100110100111001010100011000011001001111101011110110001101111001010100011100100001100010010111100110001000001000010110011111010101011110010111110101001110001001001100011111011001011100111000110101111110111001010010110011100101001101110111000101100000101001010011000100001101011001111000010110000100100111010111111000110101010100001110000110001011001000010011000010110101100001111101010110010011000110010011001100011101100100011011110101011100000011010100011001011101100000101110110100110011100101010001100001000001010101101001010101111001000010010110011110100101100100110011010101101001100010010100010100110001010111101000010010000111100101010110101111001101100011010110110110000111010100010101010011100000110100001010110101110010010100010011110101101101010011101100110100110111001000010010010110010101011110000101110100001000011010010100000101001001010110110010100100011010000100010100110101011001011000111111110100111101101001011000011011010001100000010110000101001011110101010111110100000101001011011110000101011001111100010010001011000101100010101111100101110001111010010111000001110"),
("1010011010111000101010010011010000101011100000110010001100000100101011101010100010101000100101100010011011110110001010101101010110110001100110001010100101100001101010101010111000101110101100000011001010011011101011011011110110101111100001110010100010110110101011000011110000110001110011010010101100010110001011101111111010110000111010110010110001111001001001010100011100101011010110110010010000110110001001010110101100101100111110010010111011001001101001001101000100011000010110110010101001110101000110100110100100101010111000101010000100010110001011100010011110101000101101101010010110100101101011010101011100101000000011000001110010100101001100000011001100101100000100011010111110101100001100001100111000101100010011000010010101000001001010010010111010101010000100001011000010110011101010101100011100101110110000000010110000111011001011000100111000011011001010110010100011010100001100010111000100101001100010010010001111000110001100000011001000110010011001110010111110001110000110110010011010101010100000111010000100010011101100000010111000110000001001001010111010110111101011010110001010101101000000001010100111000100101010011100111000110001101110110011000011111000101011100100001000110010000101100010110011000011101001100110010100011111100011001010110001010001001001110111011010110001101001010010100001100100101100000011101000100101110010100011000001110011101011000011010110101010100101110010111011011010101011110010010000100011000111110010100011010110001100101110010010101011101001000010010100110100101010111000100010101101011011100010110101000100001011011000110000011010011111101011001011001000101011100100111000100011001111001011000001110100000111010111011010101001000011000010110001100011001011011000100110101011101010111010100001011011001011010011101010110001010100110010111101011111101011100110011000101100010110101010101101001000101011000110010000101101010001010010010011110010101001010101110100101011100111011010100100000100101011000100111110101010101011000010110100001010101011011010001100101000101000111010110010000001001011000110001100101011010111000010110010010011101011011101110110101111100101110010111000110000001000110010111110101110111000110010011110100011001001100110011100011100100001111010101000001101001011000111101100101101101110100001101111111010001100000011011110101110111000001010111011000011001001100110100010110000000100011010101001010010001100000100010110101000001000111010111110001111101011000011111110101001001110110010111011100001001011011111000100110000001101001010110111111001101100000100001000100001111010100010110001100011101000100011010110101110010001010011000010011111101011111101111010101000001010101010001010110101101011011000101000101101110110011011000000000001001001001110010000101101111001111010110110001000101011011000000010101111010010101011000001000100101100001001000110101100011001000011000001011001001000010000000010110000100110100010010011011111001001110111011010101010100110101010101001010110001011100010110010100111101011010010110101000011101011110000000000101100110011000010111001011001101010011110100010110001111110000010111001010101001010010111001010101000011010011010001001011111001011100100000010100101000010001011001000111000101000100111111010110000010111101010110010110101001001011011011100110000010111110011000011111111101100001010000010110000001000001011001011111000101100010100011000101110011110000010110110011101001010100000111110110000010100111011000111100001001000101000110100100100100001001010100101101000101100000110011110110001101001000011000001001011001010110100110110101100010000010010111010001110101011100010111010110001100110100011000110010110101100000100111100101100001100001010100101000111001001111001111010101010111001010011000010111111101100010111101100101100100000001010101011101001000011111111111000110000001010000010110100110000100111011000000010101111001111110010110010001000001000110011101100100110110011010010100001010100101100001111010000100111000001001010111101110011001011001010111110101111010010100010111010110101001011100100011010101101000110110010110011110010001011101111001010101100110101110010011111111111"),
("0010001101001011001011111110000010101001010011100010110010111101101100001000001010101111111001101010100101001000001010101101000010100011111110111010110010001000001011100111110000101110010101000010110010100011001010110111010110001101000001110010100011011111100110000000001110101011011011010010110110010010101001001011110010110000010011101010111001000010001011001000010110101011110110001000110011111000101001010110111110100101110000110010010010111010101100000101111100101010000110111010100010110001101100000110010110110000001000011010100010000100001010011100000100101101000100110010011101011100101011000100000010101101111011101010101101101110101010000101001110101110001111111010101111001011001011110011100000110000000101000010111110011001001010101111101010100100110101111010101100011000101011011110011010110000100001110010111010000010101001010000011110101001000011101010010001000000101011110101111110110001011001101010111010100110101010000011000000110011000110000010101010101011101010000101000000101110000010111010111110101110101011011011000010100110000101101010110011111011101100011000011000101100100101011010111010010100001000000000010000101101110100011011000110100001101011110110111110101011010111000010110011111011001010110100001110101100101101010010110101111100101011110111001010110001101010000011000110110011101100000001110100101011010101000010101010011111001000101101100010100100100111000011000001111001101100001101011100101011101111100010100101100101001011000100100000011110001100110010101101101101101011000100011110101111011010011010111001110000001010000011101110101100011011011011001001000111101011101111010100101110111101000001100111001110001001011101000000100111011100100010010001001001001001110001011100101100001110000011000011101000101011011100000100101000000000101011000100001000001010010100001100110000101011010011000010100100101011010000110110110000100101100010110010111000101011100000010000100011101110010001110011000000001000110000010110110001000110101010110010011100001011100111100010100010000100110010101110011110001011000001000000110000001101110011001010010111101011110010001100101010010000110011000000100011001100000000010100101010111001010010110010010101001000010000110110101110111011101010110011110110101011111110001100100001101110010010100111101001001010101111100110110000001110011011000111101110001001100010101010101101100000111011000111001011001011001111000000010101010100111010111000011000001001101010111010110001110010011011000010100010101011100011010010101110001010011010101111000011101001010101000110101111000001101011000111011111101011101000001100101000010000000010111100110010001001101000010010101000101001111010110111000001101100010001100010101100010000011001011001010101101010111100101010100110001000011011000001010110101010100011011110101110101111010010011111110011101011110011001000101101011100000011000001001010101011000001110010101010001000011010110110001101101011100001010100101101010001010010110110001101001001101011001010101011011111001011000100011000101000100111001010101001101111110010110110000111101001010101010110110000101111101010110010110111001001111000110100010111000101100010111101000100001011110110111100101111011110111001100100110000001011001100101010110000011111011010111010101000001011100000010000101011010100100010111011100101101000110011011000101000111101110010100101110010001011110000101000100110010011111010001000111000101010101000111000101001011100111010010000111001101100000011001100101001011011110010100011010000101000001010101010100001111001100011000011001100101011111000100010101001010101011010100001101100001001011001000110101100110100110010100110110001001011110111101000101100001110111000110001101001101100001011000000101100000001110011000011010011001011100010100110101010101110011010010011110100101000100010100010101110101010100010101110100011001010110100000100101001101111001010110000000101001011100010110000101010110010010010100000100111101100010000011110101101101000100001000001011110001100001011000110101100100001000010111101101110001010101011001100110000000110100010101001001001000111011101110010101001111101111010111110101001"),
("0010101100010010001100010000010100100110011100000010100100010010001011011011011010101001000101101010110000110111101011101011110110100110011001100010101101001110101011100000001100110001011010111010110100001001001010100000010010101100111100011010111001000011101100011000000100110000011010001010111010110010001000011000110010101000110101100010100101101101001010111110110110101010010110011010111010110111001000111111111010101101111101010011000101101101001010101101000010101100010100011011000001001001101010000101001000101101111011101010110001000100101011011100001010100110101111001011000100110111101001000011110010110000000010010010110011011111001010100011000100100111010100111010011111110111001100001110000010101100111101101011000010010101101010100101001110011100010110111010111110100011101010000101110100100100110000001010101101110011101011100011011100101000010011011010010000001111101010101000101000101100010000101010110101010011001011111000100100101100111000011011000011101011001011110010111110101001000101011010011111001100101100000011111000101100000111000010111100000000101001000010000010101110010011111010100101011110101010011100000100110010011101001010011111010001101011111001110100101110101010110010110000111100001000000000000110011111110111110010010101110101101100100000010110101101111111001010110100101001001011110010010100101101111011111010100111111010101001000011011010110000001101010011001000101011001010010111101100101011001011011001110010101111101011100111101000011110001101011010000001000001101010100111010100101110110010111010110000100001001010011001001110101100010010111010101111000101001000000001001100101100010101110010100100000000101010000101011100101111000100001011000010001000101011111011000010101001010101111010001001001010101001101010001000100110110011000010110000001000101011010001110100110001110110111010111101110001101000101100010010110000110001011010111100001100101100011111010110100110000011100010100101101001100111000001000000101100001000100010011101111100101010011111111100101011111011111010101101110110001000010110100000101111010111100010100111011111001010011101111000101111100101011010111010010110101100001001110010110010000110101010011010001011101010001001001010110000111011111011000101010100000110001110110100101110110001001010111110010000101010101000110000101100100110111010100101101000101010111001100100101110010011111011000000110010001010001010000110110001101001111011001001110100001011110101001110101011000101111010110001000100100100000000000100101101001000100010100111000100001010011100110110101001011101011010110101001110101010001110001110101000001011110010101100011011001011101101001010101110000111111011000110011011001001110110110100110000001010101010110011111000101001111010000010110000111100000010110010000011001011100111001100101100000100001010100100011000101100110110110010100111101000100010100110100011101000110101010010101110000100000010111011000111001011011100101110001000101101011010101101010001001010110000010000101100011010110010000000111101101001110110110010101001111011111010110000010011001001110100110100101001101101110010110001001101001100011101000110101110110100000010110110000101101001111101011010101110001000101010110101110011001100001100110010110001000011000011000100000010000111111000011100110000010010100010110001001101101011100110011100101011100110000010011011000111001011100010100010101101000110101011000010100000001010110000000100101100001000101010111101100100001011100111011000110000100101001010011001101100101011100100100110101010111110101001110000010100001010110101010000101110101100101011000001011001001010011000010110110001001111111011000001101011001011010110100010100100010110010010111101100101001011101010101010101001111100101010111110111011101010000010011000101111110010100010110000100101001100001011110110101100100101101010111111101101001011000101101000101001100010111010101101101111101001010010010100101001100100101010111101101111101000011000110010101000100000001010010110111001000111101001100100101001111001111010111011000011001100010000010100100111000000010001100010000100001011000000010010101001000010011010100001110000"),
("1010110101111001001100011001110110101001011100000010101010100001001011111001111100100100100110111011000011000111001011110110110100011010010000100010110011001001001010100010011100100111000110100010110011101011001011000001101000101110100011111011000000110010001010111100011010101001101000110010010001111111000111000010001100101110100001111010100000000001001010011011111010101101011011101010101110111100001010110011010110110001000000010011000000100100101100000100001110101110001000100010101001011100101011011110111000100010111001010010100110101100001011001110111010101100011000101010100001010011001000011011001010010001110100111010111000110101001010011100101010101001000110000011000001001100000110011010000110101100100000110010100111111011001011000001100110101111101001100010011010101101101010000110011100101111000110001010111011000101101100011000100010101001111000010010101111101101001010000100111000101111101111110010010001000110101011111000110100101110111011011001111000110001101010001100011110101111100110111010100001100000101011101100101010101101010000100011001010101111001000111000101000101001010000000010110100011111001001001111110000110001101110001010011101111000101011001001000010101111111010010010110000010010101011011111011110110000101101001010100010011010001011001100101110101101010111111010101110000000101010011000000000101111000100000010110011010001101000100110111110110001110011110010110011111010001001001100110110110001101011111011000001011111001000100001001000110001000110101010010011111011101011001100101000101101000010001010010111011001101010010101000110110001000010001010010100011000101011001011001000110000111110101010110010101101001011101001000010110000001100001010110011011101001100001100111110101100101000011010110110011110001010010001000110101001100110110010110101101000001100011100110000101001101011001010001011100111101011000100010100100100001111110010111100101111001010110111110100101011101100011010101110100111001010010100110010101111000100000010110101000011101010010010011100101001001111111010110111110101101011000110100000101110111001110010000100001110001011001010100010100110010110011010110100010101000111011101100110101110101101100011000100111100101001100001110010100000001100011001111101000111001001010100001100110000101111011001101100001001101001001100001010100111011001100010100010110100001001000101111000101000000010000010110110110101001011101100000100110000011111100010100010011011001011100100011010110000001111100010111011010000101010111110000010100101000010100011000010111101001010100000111000101111001010111010111110101010101011010010110010101100110100110010101111111110101001010000001010100111011011111010111101001011101011110101010110101110010101010010111011101010101100010010100110101100001011101010110001000010101001110111011100101000000011101010010110100001101001001110101110110010001001000011000100101010001100100110010100101100011101100010001111101111101001111111000010110001110110101010001010100101001000010110001100101010001111100010110111110001001011011000110010100100110111011010111000101000001010010101111110101011100011101010010101110000101010000110100100101001000010000001100110101010101010001001101010101100100001110011000001100111001011001001101000101111101011011010110010010110101100001010001000110010010110101010101111111001000111101011101000101010110111111010111011011110101011010000100100101100011001100010110100010010101011001001100000101011111110011010100101010101001011000101111100110001000000110010111011100011001011100001110100101100100100000001110000101101101011010100100100100110111001101010110010001100000110111010010110101101001010111010101011010101101011000111101010101110011111110010101101101010001011100000011000101111101010110010101110100010101000101100011000100100111000111010100001010010101010011100100100101101010011001011000011100001001100000011010100101100001100000010101000100101001001111011110110100111101100001010110000110000001010001110110010101110110100110011000000100001101011101000000000101011010111011010100100100111001011110110111000110001110001111011000001010010001011011100000100110001010000101010110101010110"),
("1010111110100111101010110111010100101111001000011010010000101110001011000000001000101011001011111010110000011001101010011111110100101101111011011010110100101010001010001000110100110000001010101010101001101001001011000101110010101110100001100010001111101011001010101101100010101101110101011011000101101010001011110101000010100101011000101010110101110111001001100010111000101100110000010010010000011010001100010011000010100000010010000011000000101010001010111101110100101111000010011010111110110000101011001110011100101001100001111010111110110110001011001001100000101000101110001011000010001110001100001000000000101100110010011010101110100100001011000011100010100110011000100010100111110011001100100011110010101100010100111010001101101001101011101010100110101010100110101010000101011110101001011010010110101101000010111010111111101101101010111001001010110001110110011010110111010010001100100000000010101001001010000010110011101100101001000101001110101000100011000011000000111001001100001110110010101010000000101010110000100011001001010011010000110001111110010011000101011110001010001111100010101010100111010011000000000010101100000010110110101010000011000010011110001000001011001110100110110000111011100010110000101010101010001001101000101101110010111010110011100101101011000001000000100010101101010010101100111000001001011110100100101001111001111010101010000001101010010000010010101101111101110010110110011000101010101110111010110000111100101010110001000010001011100111010100101010001101010010101000100101001011111100011010101101011110010010101110101101101010011011101110101110111110011010110000001000101001101110101000101100101010101010111000010111101100010101011000101011011110111010111000001000101010011001001010101110010111010010110001011100001010111110010010100111100001001001110110011011001100010000000010101111101011011001110100100111001000110010100010101100100011010010111011101011101010100100001010100111000100110010110111010110101100011101101000101011110010111010100000101100001010011000100100100011101100111010000011101100001100000111000100101011001100101010111111101000001010111001111000100011101011101010110101000110000110011111011110011011110001010010101110111001001010100101011000101100110000111010000001101101101011001110100000101111111110010011000100001111101001001110100010101101110111010011000010011001101011001111111000101110010010011010110110110101101100000011100000101001101010011011000001010100101010001100001000101010010100101011000100101010101100011001011100100001011100010011001000010111001100100001101110101101001001011010100111000110001100000001010010101101000010100010111011011000101010000110100110101011111001110010101011101001001000110110010100100011111000011011000010010111101011001111011100101010100101011011000011010101000111111011111000110010000110011010010100110111101100000100111010110000111100010010101010100000001011000101110110101100000010101010110001000011101001010011000000101100000000110010101010011000101011001001111110101100001001100010110110001000001001010110111110100100010110000011000101000101101001110100111010100101100010011011000011000000101000010101110110011001000110011010111110110000000111101000000100001100100010101010100011011111101001011110100100101110000010001010100000111110001100011000010000110001101101000011000010111000101100001001001110101100001110111010111000001011001011101111110000110000010010110011000001001001001010110111011110110000001011111001110000111111001011010001010100110000101110010010110111100101001100001101000100110000001111000011001010010110000010110110001110101111001110011010100101000011001011100100001100101010101011011010101001000110001011001111000010101010101111010010111111100100001100010010101000110001110001010010011010001101101010011000001100110000101011111010101110110101001011011100110110101100110100101010111100010011001011100101111110101011110011111011000000001001001000110110010000101110110010101011000001101000001100010010000010101110001011000010111001011001101011011111110100110000110001011010101011101100001010001111101100101110001111010010110010001111001011000101101110101001101001110010000111101011"),
("0001101010000100101010011011011110110001100010100010011110000010101010000100100100101010101000000010111000111101001000010100010110101100001111110011000000101010001010011011011000101110110100101011000001010111101011010101001010101111100010111010110000111111101011111011010000101110100101100010010100101010101100011100000110100111000011001010011000110111001011110000000100101110110110111010010100110001001100001111101110011100011000100011000011010111001011000000100010101011010001000010111000100010101010001101010000100110111010101010000101001010101100010000010010110010010110110010110000101011001000000001001000101101110011011010000100110001101011011000010010101001011000001011000000101100001100010111001000110001110000111011000001000101001010100111111000101011101000111010110101110111001100000011000000100110011011111010110101101001001010110001010110101011110111100010111111100011001100001001100110101000000010010011000011010010101001011110111010100011001101100010010110000011001011001101010010101110100000111010101110001000101010011010111100100100000110000010111001100101001011100100111110110010010101001010100110111001001011001000001110101110110001101010011111001011001010010111001000101100011001000010101110000011101011100000001110101101111000101010011011000000001011101100100010101100101001111010110101111010101000111010011110101000111111000001111101000011001011011001111010101001101100001011000010101000001001001101100000101011011100101010110111001101101000010110111000101101001110000011000100011101001100010000100000101010010111011010011101010100001100000000010010110000100111100010100000111100101100001100110100100010001111110010101111011100101011100100000110101010001101000010100010001100001011001110100010101011100010011010101001111111001100011001000010101101001010100010101001011010001000100000111010101010110110010010110001101111101011000101001000100110110011011010100111110000001100010111100000101101011101010010110000011010001100000111111100011111010101001010111110101010001010100111101000100001111010001010111101010111001100100111110010100000110000010010110111001011101011110110011100101110100111110011000001100100101100011101011110101010110100001011000110111010001011001100011110101100001011110010110011110011101011010100110110101000010010010010011101111011101001001110010100101000000111110010100111010111001010100001000110101111101000001010111000111000101011010101011010101101100111001010101101011100101010100101100110110000011101011010110110111101101010111010111010101001001111100011000011100000001100011101101010101110011011011001111001111110101011000111101100101101000001010010100101101100001001111111100100101111001010000010011111010101101011101001111000110000000010111010110010011110101100010110100010101011011101111010110111000011101010110110011010100110101101011010100001001011101011001000000010101111100010111010000000011000001000100110000000101101110001100010111111101101001001110010100110100111100000000011001000000100001010011010110110101111100111110010101001011000001001110011001110101111011100011001110110100110101011110110111110110000110100101011000011111001101001010111101100110000010111001010100101110110001011011011011010101011100110101010100010101111001001110100001000110000111011001010110110100110001000011001011000110001100111010001010011111101101100001101010110101111001100010001111001011110001011100001110010100101100111100010110110111100001100000110111000100110101010000001100000011000101001000111101010101010000101100010100001000011001010011100100110101101111100101001100010110100100111100111000110101000010110100010000001000110001000001101001010110000111111111011000010101111101011000010100100011000001111101010100101000110001001011011110100110000011000010010110001110100001011111111011010101111100100111010110100000100101011011000001000101101011010111010100110001010000100000010000110101111101000010010100100110010101011101000101010110000001001001011001001010010001000100000000110110000001100110010111001010000001000000111101110101001011001000010111011000001101011000101110110100011001011110001110110011101001011001100000010110001011100011010011010101100"),
("1010100101101000101000001001001000101001000001101010001001001110101011000010101100101100101001010010110110100001101011101100111100101110001100011010101001111100001011100110011010101101010010010010101010110001101100001001000010101011101000010010111001101011101001001000111110101100110010001011000100011111101000010100000100101110001101100010111001011011101010101110111000010111111100010011000101000011101000001110001110100001000011111010111000110000101011011101011010101010111100011011000000001010101100000010000010101101011011110010111111011010101011101000011100101110010000111010110100011001101011111010100100101110100011110010111111000011001011100101110000101001101001111010110100100000001100011011110010101101000101101010100000100100101100010101010010011011101000110010110100011000001011100111010010101000111011110010110100101111101011010000010110101100010111000000111011010001001000100110111110101101011000100011000000000101101011110101011000101100101001111011000011011111101010111100011100101100110011000011000001100001101011111000010010010000101001110010101011101100001011000011011110101001111001011011001000110110101011000110110000100101111010101010110010100010101100000100100000100100010110110010100011010111101011011010111000101111001001101011000011100000001010010001000010101001100101101010010110010100101100000001101100110000001110110010101010001000001010011000000110110001110011001010111100111011101010111011111110110000001111010010100000001110101000111111010000100010001101110011000100110000001011110000001100101110101100000010110011110111101010000110011110101101111011101010101110001011101011111001110100101010110100100011000010101111101001100111010100101010100111000010010011010111101001000101101110100110101000010011000000111101001011010010100100101110011111000010011111100111100110111001000100101111111101011010111001010111001010001111001000101000010101000010110011000100101001000110001010101111010001101010100000100111101010011011100110101110000010001010100101101000001001010001100100110000011000010011000011010111101011000000101100101100000101010010100010010010001011101001011000100010011101110011000100011000101001011111000100100111110001010001110111000111001011101100011010101110010000111011000000001110001001101010110100100111011111000010100001101010001010010101010010101101101011010001001101111111001011111111101110101101011100010010110001110000001010001011101000110000101101010010101001010101001011101010101000101111100111100010111110111010101100001111011100101111011101100010100001000001001100001110111100100111110101000010000000101000101011001101110000110010000000110010101111101000101001001110110010100000011101110011000010010111101011100101110010100000001111010010110111111111001011001001011010101100001010101011000010011111101011101101011010101100101011010010001101110011101011000001001110110000001000010010011101101110001100011110100100110000000001100001101010001111001011110010001100100110101110000010011101101100001100010010101000101000011010001010110100101100001011011010100000011011001101010010111100110100101100000100110000101110101000000010111000011111101100001111110000100110111011110010100110111101001011011100101010101010101001100010111110011111001011010000000100110000100110010010101011011011101011001100011100101101000101010010110110011000001100100000010000101100000111111010111001101100101100000001110000110000001111000010010011011100001100001011011110100111011001111010110111001011001100011111110110100110111010110010110101111101101010100100010100101101001011100011000110100110001010100010000100110000101101101010011001110001101100000100001010101011101001011010010010000001001011001110110010101111011000010011000101111001001011000110001100101010010000010010101011000001001010110011100100100011101000100010010011111000001011100110111010101011100100011010000101100000101100001011011010110001000101011011000101110010101011110100110110101110110100000010111100001000101011010000001010100100101101111010110010101001001011101000001100110001011001110011000001101111001011011010001000110001100101100010110100010011001010111110001010100100111101110010000100000110"),
("1010111110111100001010001010010110110000111111111010100000000101101011001010011110101010101101010010100010000011101011110010001110110000010101010010100111110111001100011100101100110001010111000010110010000010001010001100110100100110100010000010100111101110100111111111101110101100110110001010111011101100101010011010101000110001100010010010110101111001101011000001001010110000010100101010110011011000101011101011001100101110100011010011000011110011101011101010011100110000011011100010110000100111101100010010010110101100101101101001111100101110101001000111011100101010110011100010111100101100100000100010000000110000001111000010110111000000001011001010100010101101110100111010110001000010101001011101010010100111000110000010010101000001101011100110111100101111000101101010101000011101101100001001101010101110001001001010110000100001001011001110000010101100011010100011000100101010101100010010011000101100110001010011000100101000001011100100111110101010100100010010111110001010001011101011110110110000000010011010101111010001101011011000001110101111101011101010110001100010101010110111011000100110100101010010110100111101101011100100101000101110100110010011000000101001101011010001110010101110011010001010110000101100001001000010110110100010000001011001100110100100001100001101000110011100010111011010111001000110101100001111000100101101000010100010101000000111001011110001111010101100001001101010101100110000001010101111111000101101011001111010100100011100001001110001011000101100101000010010111111010101101011000000010000101010111100110010010110101011101100001000001000101010011001101010010100000011001011000100100010110000111100110010100110000010101010001111011110110000010010110010110110110010001011001010010110101101000000100011000000100001101001101001011000100110000010011010100001010000001001001111100110100101001101011010100011010001001011101011101010101010000011000011000000110100001001000001011010101100000010110010100011101101101010000110001110101000101010101010111001011001001011100010111000100101100011101010110010100000000101010001000110110000000010000010111101110100101011010101000110100000111010001011000000111111101001101100001100101110110011011010110000111111001000011011000000101000101111000010100101000100100110011011110000110001100010010011000001011010001011010001111100101110000010110011000000011010001011000001100010100010111111100011000010000011001100000011101000110000001011110010111101101111101011111111010010110000111010100011000111100100101010100110110110101100101010111011000011011101101100001111000100011101110011001010111001100001001011100000001110101100100100111011000001110111101011100011100110101011100010101010111011110110100111011010011100100011010001011001000000000110101011101010010110110001111101001010111111111011101000001010001110101101011110101010100010011001101011100100000110100100000110100011000000101111001011010101111000110000001010111011000011010100001100010001101000110000011101110010010011011000001100010011100010110001000101101011000101001100001010110010110110110000001000011010011111111000101010001000010100101001100111001010010101000011000111111111011100000010010010001010111001011010101011100001010100101111001010000010100111011110101011011010110110101111000010100001111110001111001011110110110000110000110100011011000010000011001010010000000110101101101110010010010010111101101001011111111100101000000100000010111010111111101000110110110010101011010001110010111111001010101010011111001010011100001110101010111001100101001011100000000010101101011111100010001110110000001100000000100100101010011000111011000101000001101011111100011000101000000110111010110110000011001010110011111000101001011011000010110001110010001100001001011100110001010110011010100111010101001011100110011100101110101101001010010000000100001100000010111100101011110000100010101111010101101011100101110100101001000000001011000101110001101100000001011010110000001000011010111010101011001011111110100110100001000101101010110000011000001010011110111110101000011101011010110001110111101010100000101010101101100001011001101100101110101001111001000100101111000011011010010011010110"),
("1010110010010010001100000110100110110000001100111010111100110110101011110001110110101000001010111011000101000100001011001001001000101110111101111010100100100001101010111001100100101001100110101010010101111100001100010011010010110000011001111011000001101100000101100101110100101011001000011010101110011101001010000100100110101100011010000001101100011011101010100110101000101100101111010010111111011110101010000001110000101010001100011010011100100010101011011100100000101110101011100010010100111101101010011010011010101101101001001010111101101000101011001111011010101001100001110011000000011100001010011011011000100110001110100010000100111101001000101110111110101111111101100011000101001101001011111100101010101110011001001001111100011011001010110100101110100101000111011010111101010010001001110111010010101110110010010010101001100111001011111011001100101111010111010011000001000001101010011110110010100111111000011010101000011010101011010110100100101101011101001010111101100111001001001000100100011100001000111011000010010111100111010011101110110000001010010010110110111001000111111101111110101110001001100010111001001010001010111100000110101001101101110010111110101011101001101001110100110001000110001001010011111001101010011001100110101101111111101010100111101110101011101111101010100000100010100010101110100111101100000110101000110000110001010001111111101001101011101110000000101100000001101011000101100010001100001000010110110000101100110010111011001100001011111100011010101100100001000011000101000011101011010001001110110000011011101010110011011010101100001110011000101110000011000010111110100100001010101001110010011110101001101010110110001000001001010001000010101111010100100010010000111001101001011001011010101011101000111010101010010010001010110100110010101001111000010001100100111110101011000000001000101110001111101010101110110010101011001100001100101101010000110011000001010100101011000010110110110010001010101010101000001100001100000010010010101111111110101010100001011010101010100100010000110001100010100010001101001001001011010100110100101110110000111010010110000100101011111111001100110000110111101010111101011000001011110011010000101000010111001011001000010111101011100011011000101011101011101010110111100000101010011110011100110000011101010010110110000111001000001100100010101101100110000011000000001010001000111100001100011110011111001010100001100011101011110110010100101110110100010010110010010000101100100101011010110000110100100011000000000111001011000101111110110010011101000001101001110111101011010110011000101010010001010010100010011110001011001000111110101100000000110010011001000001001010100011001010101000010010110010011000011011101011011000111010100000011011101010111001010111001010000011100000101001010110001010101010001010101011101010000010100110001101111010101010011011001010110010101100101011101101101010111111001111001011001001000000110000100010101011000011100010101011000111000000101111000111000010110101001110001011101100000010101111100111011010111111010101001011011111001100101100110100100010101110110000001011111000011100101101010100101010101010000011101011001111001100101101101011000001110001100001101100010001111010101100001111010010110111000001001001101100100110101101000001011010101111010000001011001101000010101001100001011010100011011000101001100000110010101100011110110010110000111110101011100001011010101111100100110010111010100010101011110010001000100100100111100010111111010100001011110000011010101110010101001010011111001010001100010000101000001100010010000010110100100010001010001000000100101100000111110010111001100001101011011010101000101100111000110010111101001010001011101101010010101101001111111010100000000010101011010011000100101101010100000011000010001001000111100011010010101001100000011010010111010001101000110011011100110000011100100010110000100111001010000101110100100011110010001010110101000110001011100001110100100011100000010010100001000110001010010111101100101110010100001010111010011011101010111000100000100000100010010010101011110111001011101000110000110000111100100010110111111000001011100001001100101110111101111011000000011001"),
("0010010111101100001011011101001100101001100101111010101011111111101011101011100100101011011110110010110000011100001100001001011010101111011001111010110001010000101010100101011000110001001001011010010111010011001010100110100100101110000111010010111100010110001011110110111000100001010000100010000110001001001001110011011010100100010111101010000100110110101011101000000000100110110010101010111011111010101011010010110110101101010010101010101011011110101100001110001110101111100000101010111001001000000111101110110100101001101111111011000000010010101011010101000010101100111011110011000010100110101011011110111110100000011100010010110110100100101001010001000100110000000011000010011111100010001010101010001110101010001100101010110001110110101010001100001010100100011001000010010101110110001011011111110000101011010111000010111011001010001010110001011000110000001100001010111100101000001011110011011010100000111010001011000010010010101011001111110010101001101100010010110001101011001001010001100010100001100011111010010001100111001011011110111010110000110110010010100110000110001100010100001100110000010011110010101000001101001010110100010110101110110001011010111000000011101010000100001000110000010000111010010110100111101011111111101100101010000000000010011000110010101010100111110000100100101011101011000100000000101100001111101000100101100101111011000011000010001011100001100100101100001010001010110010111000101010011011100100101100100101000010100001011101001011001100011100110000001001010010001111001011001100101110101010100000010011110011000100011111101010101101101010101100001110110010111110000010101010001110111110101000111010100010100001011111101100010100011110110001000010010010101001111000101011110010100110101100000100010010101110011110001011111011001100101100000110010011000100010000001100100001110110101111011011001011000111010011001011110000000010101001010010010010101111101110101011011101110010110010000010000010110110010000101011000100011010101011011101000010010100100110001100001111100000101101101101110010111111101000101011010001011110101011100100011011000111010001101010100110001110101011111100001010110010001110001011110000001000110000000110110010101001100011001010101000111110110001111101111010101101010101001011010100000000110000011100110011000010101000001011100101101100110000100001100010110010101000101001100001011000110000001011111010000011001010101010110010110100101110001110011011000011100101001010111101100000100111000100001011000010010111101010000001011100101001101110010010000100110111001011110110111000101110111011001010110111111101101001001110100000000100100011101010110001110110101010011110111110101100000011001010100001101100001010001001100000101000110011110010110100011110101010000011101000100110011001101010111010011001101100000001111000101110111010001010101010001000001100011011010010101110000110011011000001100011001011101110010100100110011101110010110011001001101100001001100100101100110010101011000000011000001010011011001100100100110110110010101101101011101011011000001010101000111100011010100110011000001100011101001010101110100111001010111011011101001000100001110110100001111101011010100010110001101010110010111000101010110011011010110100011111001010100010101100101110100001010010101010010011101011001110000100101110000111011011000001000100001001101110101010101100110000110010101001010101101011011111001000011010000111001010110000101000101010000101110110110000011010001010110100101001001011011010101000100100101001011010100101010001001100001010011110011100100111110011001001100010001010110101011000100100000111011010110010010100001000001110010010100111111011111010110010001011001001110011001100100011100010000010011111010000001001110000101010110000111010110010110001010111001000110101010010011110000101110010111010110000001011011000111000101001010000010010110001000001001011010100101010001101001101000010110001010000101011110000100010101100111001101010111001011000001011101111100110100100100011011011000000011000001011100001001100101111010110100011000010001000101011011110001010101110001011010010010001110000001010000100001010101010101111101011000000100011"),
("1011000010111111001011100001111110101111010010010010110001000111001011001000111110101110010110001010111010111000001011010111010110110000000011000010101110000100001100011011001100101000110000010010111111010110001010000101001100101100110010010010111101100101101011011101011110101011000100101010110110101010001100001001011010110000100110000010110101000001101100010000000010101010011001000010011111111010101011011100011100010111101010011010100001001001001001011101010110101011001001001010111110010010001100001101010100101110011001001001111111111110001011001101011010101111011100010011000010101110101011000010111110101000011000100011000000101101101011010001000100100100001001110010111101010100100111110110000100101110010111101011000001100000001100001011110100100100101000110010111110000101001010001100010110101001101100111011000011100101101011100010000000100111100111101010100111101110101010100000110110100011000011101010101100010100101100000000000100110000000101101010100110000000101011101110000100100100100101011011000001011010101001000000100010110000101011100010011010111011001011101001001110110000001001111010111101100100001011010110011010110000100010000010011100000101001011000100011010011111010000000011000000001011001001110010100100101000011100011010101000001111101011000101000100101100011101101010001010110000101010100001011000100111010011010010110101001110001100001000011110101001100001011011001000101101001100001101110000110000011001111010011100100010001011011000011000101000100110010011000110100110001100010000000000100100010011110011000111110100001011100001011000011111100011100010110101010011101010100101110110101111010000010010101011000111001010011100111000101110110110011010010011101001001010001110101010101000111100010010111000000111001100011011111100100110100011001010110000001011001000110000110100100100010100001010000110000111001100000110011000101111110011011010100010001111101011001001011110101100000101101010101011001101100111101010010000101000011010010010101001100100001010100000010010101010000000010010111100011100001010101011011110011010010010101011010000001010101010010101011110101101111111011011000000110110001010001100101110100010010110111010110011110000001100000001110110100111001110100011000010000110001000011111001000101010111011100010010111110110101010100111001110101100000111000010000111110111101100011000010100101111011100000010110001011100101010110111010110101010110110110001110000100011001000010010001110101110000110100010111100100000001010001111011010101000111011100010011001011000001011111000101000101111011100110010100010101000101100000101101010100001000111010010010111110000101010101101011100100101100000001010110100110000101011101100101010101100011100010010011110010011001100101100110000110000111011100001101011010001101001010111101100101101001111011011000000000000101100010100111100101001110011001010101101100010101010110111011100101111110111101010100001000101101011111111001010101001110011001010111000011010000111101010111010100101001000110011000101100000101001100000101000101110101110110010111010000000101010011110000110110000101011111010110011000101001011100101100100101000011010101010101101001101001010111110100000101011110101010010011001111111001001010000000100101110010100110010101000000110101011110111110110101000101111100010100011011101001001000000111100110000111111100010110000100100001010001100010000110000111100101010111001000111001000010100010100101001001111110010110010110011101001000110010010100101111111011010101101100111001011011011110110110000101000001010110000110100001100000101001100101111100010001010110110111100001011001001101010110000100000010010100111000111001100010011000000100101001011110010110111000101001010110101101110100100001110001010100111111101100111011110011100110000100100110010111101010000001001100110110100100010111110110010110101111111001100000100100000101110101110111011000001010011001100010110101110101100001001011010110100000100101011110000010100110000100000011010111011010111001010100111110110101110011010000011000010010001001001011010011000101011101111000010111001010110000111001111000010101100011101010010011111011110"),
("1010101111100101001010011011110010110000001100011010100110111000001011110010101110100001100000101011000011001101101011000100101010101111001010011010010011111001101010001010011110100100000100000010000011111001101100000000010010110001000000110010110010011010001100001001011110110000000001110010100111011100101011111100011000101100010001101010101101011010101011011100100100101100001000111011000100111100001100001100000100101101011011100010111100110110101100001001100000110000101110001010110010100100100101011011101100101101001100111010100111000100101010010011000100101010111101110011000000000111001011011110001010101111000010100010110100111011101011111101010100101111011101100011000011101110001001001010111110010111010100111010111101000111001001100101110000101010000000000010111000000111001011101100000010011110011101100010000110100000001010010001011110101001101100010010101110101101101001110101001010101110111011100011000011001110101011001001101110101100011111000010011111000100101011001100110000101010001100111010110010101101101011010110110110101010011111111010100101011011101011100011010100101101101001000011000010001111101011100111100100110000001010110010100001001000101000011000101010101001111100000010111111101110001001111111111000101111111110000011000001000011001001010111001000101000011101001010001010100110001011000001010100101010011100000010110110100100101011111101011100010101010100100010111011000010100110001101011000101000011100110010101001000011101011100110101110100011000010100010101110111101101010110001101110101000000100001001101000001111101000010110111010101100111011000010111111110100100110100000010010110000111110110010100010111101101011110101000110100011111010011011000011100110101010011000001100101000111010000010110101010111001011101111001000101000000101000010111010010110001100001001000010100011100010111011000011001001001011110101010110101000101010111010100110011011001010010111010000101000011110011011000111011100101011001101011110110001110001011010111111100001101011000010111100110001110110110010110011001101001010001101001110101101111011011010111000100000101100000100010000011101100011000011000000010001101001010011100110101011101000101010100001001110101010011000000100101000001100110010011110100001001011100110110100101011111110110011000010111100001011010000101000101100101110111010111000011101001010000011001010101000100011101010100011001010001010010110010010101010010011110011000000011011001011100011101100101000110010110010100100000111101100001001000000011110101100000011000001110010001010101100001000100101101111111001101011110101001010001001010010110001110001001011000101101101001011111000011110101111100101010011000001100001001100011111110010100100110101110010111010001100001010011001110100101101011011010010110000011011101001000110111100110000110010111010111011011011001010001001001010101001010100100010110111100010101010010011001100101001000111100010010010100110001010001011011000110001001010001011000000100011001011010010000100101011111110000010011001011110101011011100101000101101101010010010100000000110101011111100101100110000010011111010110110100110101011100100011100101101010111001010110101001010001001011111011010101011101110001010100000111111000101000111101110010111110000010010001110100010101010111111101010101011001111000010110000101001001011000110101100101110011000011010110111111110001011010110011110101110100001001010100100000010001100010100101110110001100001110010110111000101101011000001000000110001100111111010111011110111101011110111011010101001100110001010110110010100101011001101100100100001001110101010010000101010001011101001010100101111001101000010010000000100001100001111011000110001000100010010111000100001001011001000001110101010000101010010110001000100101011011100101110101101011100010010011000011100001011110001001110101011001000011010111100100011101010111000101110100110010000001011000010011000101010111111100000100001000011100010111010100010101010000101001000110001110110000010110010110101001001000000110000100111101111101010000010010010001011000001111100101110000011010011000010000001101001101011111010101101110111001010010011011111"),
("1011000010010011001011101000000000101001111011111010000000110100101011000111011110101010101011110010111111110010101010001001111000101001110110000010110101011101001010111111000000101111100001110011001001000111000111000111011100100101001110101011000110111011001011011110010000101100001100101010000011101011001100000111101100100101110111110010011110010100001010110010101100011001011110011010101000011000001011000001010000110001110101100010111100011001001100001110010100101100011011101010110010100011101100001110000110100001001110001010110000101010101100000110011110101110101010101010110111010001001010111110110010110001000011110011000010000110001010010010101000110000100000100010100000011111001011001110000000101110110101101010110000011001001010000111011000101011011011111010101111011101001010110001100010110000110001101010100111001001101011100110000000101110101110001010100110101101001011000100001110101111011101000010110111100000101010011111011100110000001010000010111101000100101011110100101000101001110010000010111110000100001011010100101110110001111000111010110001110001001011011010111010110000010110111010111100000011001011011101010010011001000000111010110010010100001100010000001100101011101000001010100001111100001011000100101110101111110110000001111110111110001011111011001100100100011001111001011100011001001011110111010100101110110111100010110000001101001100001000010000101010100110011011001100101000101011110101100000110001010101001010110110111101100111110010101000100100001000000010011101101001101010000010000000101101011010110010110010110011101100001101100100100110111001001010010111000001001100001010000000110000100010001010011011010010001011001001111000110000100001101010111011110101001100000011011000101011001101011010110111100110001100010010110010011100101010111010110101100011101001000100100100101001100011010010110010001100101011000001100110101110001011101010010001011010101011001110111000101100111101011010101010011110001011010010111110110000101000101010110010110110101011111111110110101000110010110001101000111100001001000001000010100011110111111011000110011000101100010000111100110000011100110010011001011110101010110111110010100000001101111010101010001001101100011001000100101101101101100010000100100011101001000011000000101100111110100011000111101110001100000000101000101111011001000011000001011010001001101000101010011000100010011010110110101000001010111010001000110000001010110010110100101011101010010010001110101111110101000010100001111110001011111000110110101001011111100010111001100001001011110000001110101100011010000010101011100111101010100011001110100110111111000010011100110001001010110110010000010110000111101010011101101101001011000101100110101000100001010010011100010011101001000100101100110001110101001001110111011111001011010010110000110001110000010010111110011000001010011111001100100001011010011010010010001011001100000101101100011001010011100010110010011010101011011101011100110010001010101001100111000001101010110011001000101011011011110010100101000111101001000001001100100100011000011010110111000100001010001100000000101101001111011010010001000010000011110111011110100101100000100010111100111001101011101010011100100010001011100010100010110001101010100101101000101101100110101010111011010111001010001000011100110000101100010010010000001101001011000101010000110001001000000010101111101011000111010100111110101111111111010010110111111000001100001010100110101111110010010011000101110011001010001100111110110000100011110010101000010110101011001100100000110001000011011010110011011011001011001011011010100100010000001010101100010011101000100101110110110000011110111010111110110101101100000000001000101000101110100010110111001110101011101100001000101110100010100010001000001001001010001001010100101110101010100011000100111111101011011110000110101001110111000010100101000001101010010111110010100101111010010010000011101110101001101101110000101011010010000010110011101100101010110010010010101100010001111011000111000101000111100001001010101100011011011010100011000110101010011101110100101100111000000011000100010111001100000100110110101110001011011011000111010001"),
("1010110011101110001011110110100010101110001111100010101010011110101011000110100100110000100001011010101100101111101011000001011100110000001111010010011010000100101011101101110100100101100010010011000101101010101001010010001100101010000100100010101110010101001010110001010000101000101001100010110111011000101100010110110000101101010011110010110100100111001011100001001010101101100011100010010100110111101001100001010000101010010010011010011100000001001100011101010010100110000000111010110010001100101011111110100000101111011010111010000010001011001010101100000110100001011100000010111010000111001011111011000100101000000111010010110001010000001001000010010000110000011011011010110001011101001011011100111010101101101100011011000000111110101100000010101010101111011000010011000100101010101100010000000110110001000010000010011001101010101011101011000010011011110101010001010001010101101011111001000000101011010000110010011111011010001001110110010010101111010001011010110111101010101010010011001010110000000001011010101110100010001011000010010110100001101010101011000010100100101010001101110110011011001110000010111100100001101011000001100000101011001010010010110001000111001100000000000110100100000001100010110101001010101011111101110100101110001110100010110011001111101010001001110100110000000001000010111000101101101010100100100100101000101100000010111101100010101100000110000110100110001101001011000010011100101011010110000010101100110100010010010011000101101011000011010010100101001001010001110110101010101001001010101100101000101100011010010101001001101100001011010010101110001101110010001100001001001011000011111010011101100111101011000100000001001011101100000110101111101001100011001000111100101100011001100110110001011101110010110001011110101011001001001110110000100101010010101001000010101010100000100010101000101001001011000010000010001100000001111010101100101000111010110000101000001011110100110110101011111110000010101001010000101010111010000110101110011101010010111110100010001011111011001000101101100111111010110101000000001010100011101110101101100000101010111100101100001000101001110010101011010110100010100111001000001100000110011010101001110000001010101000010110101011000000111110010110100010011010101100001101101011001011011110101101111101001010101001101100101011100010111000101100100011000010110011100010001011101010100110101111110101011010111110010010101000011011010110100101000001100010111010010001101011100001111100101111000111111010110111001000001001010100000100101101101011100010101001101001001010011010010000010110101101110011000001111101101010001001000000101001011111111010001100101110001010011101110100101111101000001010100000110011001100011110100110101100011010100010101001011110101010001101000110101100101100111011000101011001101010100101100010101101000001110010010101000010101010111111110110101000000000111010000110110011101001100011100100100111111000000011000001001110001001100000011100101101111101111010110001001101101010110110101110101110001000000011000101111101001001101000010010100100010110110011000000000110100110111100100000110001001001100010111000101110101011011001000100100010001011010010101000111011101100000100010000110000111101111010110100110001101100000011101000101101110000000011000000000010001011100110100100100111001101101010110110111011001001001000100100101011101011010010001111110111101011111001010110100000100011001010111010111110101001100000001010001011110011000010111011111000001000100100011100101000010101010010101101000010101010001101011100110001000110100010100101001000101100001001011010110000100011111010110001000001001011001000110100101100100100000011000010111010101001010101010100101110010111110010110010001000001100001111010110110000001001000010111111101111101011101100110110010011011011101010111000001000101001011001111110100000101100100010110110000100101001001010111010101001100001000010111101000001001010111111000100101110111001101011000011001010001000111110000100101110110110000001101000100011101010101010010000101100100011000010110000101110000111111111100000101110100011110011000110000011001000000111000010101100011100101010100010000000"),
("1011000111111001001100011010000100100100111011101011001000000111001011001100011000101000001100011010001110111101101011010101001010100000100111000010111101100101000111111001000010101110010001010011001011010011001011011101101010101111001110101011000110011110101010001010110000110011010101111010000101010100101100011000101100110000010111011010111100011011101011100011110000110000100111101010110100110100001011001001111110100010111011001010000011100101101000101101111010101011011000101010110100011010101100010000101000100111000010000011000001110000101100001010111110110001100100111010011010101111101010111000010100101111010100100010011001111100101010010001001100101001101001110010111010100111101011011000111100110000001001111010011000111010001011110100111000011100100111101010111111110010101001100010001010101010011110001011000000111101001010101100101000101100100101110010111100111000101011101000101110101101110010100010101010110010101010011111000110101101111001110010101011111111001010010100010010100011011001010010010101110101101000111111111100100010011110111010101000101001001010011010010000101110110011010010111101000001101100010001010010101011010010100010011000111100001011000110000010101010001111110010010110111001101011111100011110101111111010011010010110010111001100000100011100110010111100100010110010011001101011010011100000101010010111001011000100001110101001110010101010101100001001100010101110110010101011111011000100101111111101111010100011101100101011000100000000100110001011110010011011000011101010000110010000101100001100100010001011011111001010010110011010101010100110100011000011111101000110011100101100101011101110111010011010101000001010010101100110101111000101010011000001111110001011011001011110101101111011101010101110000001001100000010001110011101000000011010010011101001101001000111101010101111001011101010111001000011101011001100111100101100001001000010111101110100001011110000001000101101010110110010110101101110001001100011001100101011000110010010000001011000001001101011110110101000111001111010110001101001101010000110010100110000011001111001110111101100001010011011001010101010100010000010001011110011001011010010000100011101010101000010101111110011101010011011110010101100111100110010111111000000101001001101100110101010101010100011000001001001100111100011110100100011100111111010011001110000101010111100000000101110000100010011000100110111001011100100010010100100011011011010111001101110101011001111111010101100000011010010000010001010001100010100100110100010100011110010100101011000001010001000000000101100110000100010110000111001001001111110010000110001001011011010100101100101001011111110100100101000011100110010110010111001101100010001010010101100001000101011000001110010001100000101110100110011001011001010100100000100001011001000100000110000111000110010010011000000001011010111010110101101010011000010111111010111001100000010010100100101100100000011000001001110001010000001110110101001110111111011000001010000101000110110011010100101010100100010110110010011101010110100100000101101011000011010010111111100001100011000000000110000010111001010011111101010101011011011000110101011010011100010011111100101001011100001110110101111100110001010001111100110101010000011110010110001010001110010100001000010101011010000101100101101110010100011000011100000001011110100100110101100000101011010010010001010101010001111111010100111010000110010100010101100101011010001111100110000000010010010100010101101001001110011100000101110111101101010111000010101001011100001111100110001011000110010110001001111101011001101101010100110111101010010111110000110101010101000011010101110100111010010100111001100001011111100111000100111101000010010110011000000101001111010000100101001011000011010010010110001101011011110100110100010011011110010110101010101101011010000100000101001101001100010101011101011101010111001100010110010101100001010111001100100001100011111011110011000000101001011000010101100001100000111100110101110001011100011000000010100001011101001111110101000101110100010110110110111001011010010101010101100000111011010011101100001001011000000111100101100101100011010111110100011")
 );

 TYPE fixed_point_array IS ARRAY (natural RANGE <>) OF std_logic_vector(15 downto 0);                                  
 constant bias_array : fixed_point_array(0 to 15):=  (
 "0010001101001100","0010110110001101","0010110011000001","1010001100100001","0010101001110110","0010110100010100","0010010111011100","0010100000010011","0010100100111001","1010100010001010","1001110110000010","0010101110011001","0010101011111010","0010011101001110","1010101001001000","0010010000111001"
);

 signal  reg_Layer1out : fixed_point_array(0 to 15);
 signal weighted_sum_array : fixed_point_array(0 to 15);
 
 
 
begin

  gen_neurons1: for i in 0 to 7 generate
    N: Neu_Ron generic map (N => 256) 
    port map(
      clk => clk,
      inputs => layer1_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer1out(i)
    );
  end generate;
  
    gen_neurons2: for i in 8 to 15 generate
    N: Neu_Ron generic map (N => 256) 
    port map(
      clk => clk,
      inputs => layer1_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer1out(i)
    );
  end generate;

  -- Update output
  process(clk)
  begin
    if rising_edge(clk) then
      Layer1_output <=   reg_Layer1out(0)  & reg_Layer1out(1)  & reg_Layer1out(2)  & reg_Layer1out(3)  & reg_Layer1out(4)  & reg_Layer1out(5)  & reg_Layer1out(6)  & reg_Layer1out(7)  & reg_Layer1out(8) & reg_Layer1out(9)& reg_Layer1out(10) & reg_Layer1out(11) & reg_Layer1out(12) & reg_Layer1out(13) 
                       & reg_Layer1out(14) & reg_Layer1out(15);   
     end if;
  end process;

end architecture structure ;

