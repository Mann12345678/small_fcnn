library ieee;
use ieee.std_logic_1164.all;

entity layer3 is
port ( 
       clk : in std_logic;
       Layer3_input : in std_logic_vector(511 downto 0);
       Layer3_output : out std_logic_vector(511 downto 0)
       );
end entity;
    
architecture structure of layer3 is 

component Neu_Ron is 
generic( N : integer := 4);
port ( clk : in std_logic; 
       inputs : in std_logic_vector( ((N*16)-1) downto 0);
       weights : in std_logic_vector( ((N*16)-1) downto 0);
       Bias : in std_logic_vector(15 downto 0);
       weighted_sum : out std_logic_vector(15 downto 0);
       neuron_output :out  std_logic_vector(15 downto 0)
      );
end component;

type weight_array is array (0 to 31) of std_logic_vector(511 downto 0);
signal weight : weight_array := (
("00110011000101010010000100100011101011101101010010110000010111011010001101010000001101001011010010110010000011001010101110001111101100100111101110110001111100011011000011101000001100000000100010101011111011000011010101011110001011110100011110101110011111000010101011010010001010100111001100011100010011110001110001111101001001110101010100110100111111011011000001110101101100000000110010110011001101010011001001011111001100011110000110100010101100000011010000101010101100101010001000110000110000000011000000001101"),
("10110100010011010011000000101001001101010111110000110011111111010010111001110001001011101000001110110001110000011011001001011110001011000101011100110100001000001011000011111110101100100001010000110000001100101010110000101110101010000100100100110001101110100011001100001010001101001001010010110100111000011010010101000101101011010100100000101001010100011010111011001100101100101011101000110001000101001011001001010111001100100000000100101110100110000011001011010101101011010110111110101000011001101011000000000110"),
("10110100001001011011010000100111101101000110011000110000101101010011010011101000001011000001101100110001000010001011001111010010101010101100101010110100011010101011001111100011001100011100110100101001100110100010010011100110001100000010000000110011000010110011000110001100001011000001011110101001001000011011001001101110000111011100110100110001111111110010101101101111101100110001011110110000011000001010110100001001101100000111011010101101011011101010000100101100101101001001101110101110101111011011001001011101"),
("10110011111011100011010010100011001101000111000110101011001010110011000110100110101101010010110010101001101110011011000010101011001100001010100010101000100110011011001100100010101010010001010110101100111110111010110100011111101100001110010100110100101110101010010110011111101011111101000110101100111001100011010100110100001100010010000000101111110000001011000101111101101011011001101010110010110000101010100011000100001100010010001000110011011011100010110010011001101011010100110100110010001111110011001001010000"),
("10110000011100101011001111010010001011110111000000110101010000010011001010110100001100110110111100110100101110100011010000011000101010110010101010110001010100100011001011011101001010101000110110101110001111100011010000001000001010100100001000101101010100101010101101000010001100110100001000101101101110100011000100001010100111111101110000110001011000010011000100100000101011011001011110101000100111000001100110001100101011000110100110100110110100001011001111100111001011000000111010110001100110000011000111100010"),
("10101011000001101010000010101101001100000111111100101111001000010010011000100110001011001000100000110000010000011010100001110110001101010000111110101001000011011001011110011011001100110010001010110011100110010011001001010001101011111010001100110100110111100011010011001010101100010101010100110000010100110011001101000110001100101010100010110001001011101011010000010001001011001011100100110001000010010011010010110011101010110111001100110011101110100011001110010110001101000011000110101000100110111010101011010110"),
("10110001011010011010111001010010001100111100100110110010000000100001100000011110101001111001010010110010100001000011010000001011001100000100010110100110110111111011000000110000001100100100010110110100010001100010101101000011000101111110101000110101000101111010101111011001101100010111010010011111111111111010111010010110101011001100110110110100000001000011010000111001101101001110101110110000001100001010111101000010101011001111000110010010110100101010111000101110001100100011110010100011001001110011001000100101"),
("10110001011011000011001111110001101100001010110000110101100100110010101000010100001100110110110100100110000100000010110100101111001010101101101110110100010010101011000000010011001101001001100100110000010011011010111111111001001101000010110100110010010110100010010101100100001100011111011100100010111110100001101001101101001101011001011010101111011010010011000110010010001100011010001000100101000100110011001011000000001101000111101100110011011000111011001100001011101101010111100110110011101000001010101101110110"),
("10110000001101111010110101000011001010000100110010110100011100000010110010011011101000111101000000101110010010111011001011101000101011010111110000110000101110011011000100010101001100100110000010110001001101011011001111010101001010011011010110110001110101010010100010001001001101001101010110110100011110011010101000000101001101000100001010101110011000010011000101111110101011111011011100101110111011011010100000000101001100101000010010100001111111000010100000101110101100110110000100110100110100000011010001001010"),
("00110100100110001010101000100100101011000111010100101110010011010011000000110110101100010101110010110011010001000010110010111010001101010101001000110001000111001011001111001010001100111000111000110101111010111010011110000100001100010110100100110011011000000010111101011100101001001010011100110100000110101011001001000000101100101100010110100011010101010011001111000101001011111110001000101101100110000010110000011111001101001101011010110010101000000011010010001111100111010001011100110011000101011010100101100110"),
("00101110000101000011001100011111101010001000101010110010101010110011010000001101001100011110011110110101001011000010111111110010101100000101110110100110000101101001010110010001101100000110000100110011011110000011001110101101101101000000000100101110100100001010111000110000101100100010101110110000100000111011000100000100101100000100110010110011111010000011001110011110101100100110111110110000101101111011001010100101001011100011100010110100000101000011001010000100001100111111100110101000110010111010111100110110"),
("00100101001010000010011010000110001011111010100000110001110010101011010000111101101010110110001000101110001001001010011100011010001101011010011000110011101011110010101111011100000110111011100100110001011001010011000111011000101100100010100000101100101110110011010011010101101100000001010110110100000100000011000010101001001100110010110010110000100101011010100000101011001101010100000000101101000011100010100001010110001001110000100100110011010100001011010001101100101010100101111010110100000111011011010001001011"),
("00011100000100010011001101001001001011011011101100110101000000101010100010000011101100110011100110110011110100011010110101000000101000101001110100110100100101111011000110101101101100101011001010101001100000001011001000100101001011100001111000110100000110101011001101010011001101000110111100110101100111101010111000111100001011110101011100110101010010001011010000010111001011100011000010101110001111001011001100010000101100011101110010110100001110100011000111000010101011001001000100110010110101111011010001010000"),
("00110001110101001010111101110111001101001110110010101101000011101011000101101110101100000000100010110000011001111011010010100000101100010010001110110000100010010011010001101101101001001111101000110100011000011011000010010001101011000010010010011111101000110011010111001101001001111100011000100110100100110011010000101011001100101111100000110000101100101011000010111011101001010111101010110011101001111011001011010010001101001101110100110100111111011010010100111110101001000010001110100100111000110011000110110010"),
("00110001000100001010010000011101001100010101100010110011111011011010110101110100101101010101110100101000001011001011010000101001101101001001111110110011111010101011000000010111101101000110000010101100101001000010100101000100101101001001111000110001000001100011010101001111101100100101111110100111011001100010111001100101001001010010110100110011000100010001100110101101001100011111001000110101000100000011001100110110001011101100010010011000000001101010100110001111101100111001110110101110101111110010010011101010"),
("00110011110001000011000001110100001011010100011010101101101000011010111110000000001100111100000010011011101111010011001011000110001011100000001000110001110110011011001001110010101011010111010100101011101101101011001100111100101100111101001100110101010001111011000110001100001100111100010010110011101000001010110110001101101100010000110100101100000111000011000000111101001000101000010110101110011001101011001010111011001010111110010100101001111111111011000001111000001011111011011010110001100100001010111100000111"),
("10110100010111101011000100111010001100111111010100110100001001011011001000101110101100110000011010110100000100100011000110011000101100111001110100110010010111100011010011001110001011000100011000101011100011001011010001110001001011000010010110110010010101000010110110001000101101001001111010101101110001000011010100111100100110101011010000110100000110100011001011010111101011110001100100101000101000100011010110111011001100100011100010110011011110100011001111100001001100110001101010100010100110001011010000010001"),
("10110011100110111011001110001101001100001110110110110010111010010011001101111100001100100011101100110010011011010010001111010100001001101110101100110100100100110011001100001011001011110111101100110000001111000010111011111011101010000100000010110011100001010011001001100101101100010010010110110010000000111010110011011000101101000001001000101001010100110010001101000111101100000000010100110000111101111011000101101100001101001111000010110100001100100011010000011110001100110100110110110100011100101011000111010001"),
("10101100111010101010110011000010001011110010100100101000111011111010110010011001101100000100111000101111011011001011000100111011001100110110110100110010010000110011000001001101101010000110111000110010100011110010101001010001101100101010001110110010110010100011001111110111101101001101010000110000111001010011001101011100101100010010110010110100110101001011000010000100101100110001110110101100111101100010110100001101101100000011101000110101011010100011010001100000101010101011100110100100111110011011001011001011"),
("10110011010010101011000010101001001100101010000110101111110010111010111111001111101011101011001110100010010010110011001011100100001100100000010110110100110110011001110010110000101101000010011100110101011011100001110000000011101101001011100110101100001010010011000011000101101100011100100110101101001100100011001101010010101011001101111010110100001000000011010010010100101100000010101000110010101000111001110001110101001100101110101000110010110101111010110001010001001100101110001100110100110001110010101101100111"),
("00110101000100110011010001100110101000110111101100010101000011110011001100000111001100001110010000110100010001011010111010011011101001100001011100101001000110100011000001111000001011100001101100110001101000000011001001100100001101001101101000110101001001000010101000000111001100011011101110101001001110011001111111110110101011100101111010101110010000111010110110110010001100111110001000101111100100101010101000100110101101000100111000110001010111101011010101000001001001100000010010110000110110111010110010100100"),
("00110000000100101011000010000111101100110100011100110001001100000010111100100110101100110111011010100101100101000010101000001010001100111110001010101101100010101010011010000000001101000100100000110100001011111010111100110111001101001110110110101110100001000010111010011110101100110011010110101101110001010010111010111100101011010101010000110011100110010011010011000100101100011101011000101110101100111010111100011111101100011010100110110100100110100011010010011000001101000100110000101101101010110011001011011001"),
("00110100100001101011000111010100001100001011000010110010101110001010010101011001101001101000110000110100110111101010111000101000101100010010001100011001000110100011010000111100001011010001010110101100111010110011010010000011001101000111101100110001011010000010110010101011101011101110011000110011111110010011010000101100101100000110000100101000100011001011001001101001000010011100010110110100001110000010011000000101001101011001011100110100111101011011000011100000001011001101000000011110001000001011000110010111"),
("00110101001011100011010001011100001101000001111000101010010001000011000011110011101010110110010000110100111101111011000111001110101010011010011110110001000001001010011010010101001011001011110100110100010010011011001001110110101100111100101000110100111111100011000011001100001100011011010100101010110111111011000001111010101100010110011000110100110100100011010110011101000111101101111000110100100011010010110110010111101100100011011110101011110001010010101011110001001100111001000100101110010011101010110110010011"),
("00110001100000110010111110110101101101001011101000110100110000010011010110111010001011110000111000110101001100101010011000000101101100110100100100101100011000011011010011101000101100001111001000110010010111011010110111001110101100010010110110101110011110111010100101000100101100110001111010101101000011010011010000101110001100011100000100101101010110000011010111001001001100100011100100110011001010011010000111111100001010000000001110110001000001000010110011010011001010001011101110110100010111000011000101111100"),
("00110011010000101011010000011000001000111101111100100000001100011010111001110111101100011110110110101001111110101010100001101100001100011110111100101001011101100010111011100110001011101100101100110001010010100011010000000101001100100011101000110011100001010010111000100000000110111011010000110001110000100010010111101001101101000001111000110100000001100010110001100101001011111111100110110010010001100010111101111101001100101001101000101100100000001001111001010101001100101011001010101000111100001011010001010011"),
("00110011001010011010111010101101101001100011000000110101010101011010110110111111101010100001110000110011001010111011000111000101101100010010110000101000011001100010111101001101001101000001101000110000111000101011001111010010001011010110001100110011011110000010111110010011101010011001000110110100010010010011001000001000001001010111100100110100111000000010111111101110001011100111000000110001101110110011010101101011100110010100010110100101100111101011000000001001001001111111111110110000101110110011011000100001"),
("00110000001000010010010100110111001011100101110010110000001001000010101101010101001100001101110000100110000010001010101010101000101011001000001010010100000000110011010100110100101101000001111100101000011111000011000010101011001000101100010110100101110100011011001000011011001100100111111000101111101001111011000110001101101100100100000010110001111111101011001100011010001100111100100100101100100001100011010100101100101011110011001000110101100001010011010011000100001010000100101010110001110001110010100110001000"),
("10110000001001100011000111111110101011011101110110110000011111111011001100001100001101010010000110110011001001111010011011111110001001010111000010110011111000111001110010011100101100111011010100101100101110011011001011001001101101000110100100101001011100101010100001111011101011100111111100110100100110111010001100001010101011010001010110101110000110010010010010000110101100111010110000101010111100001010110111011100101001110010101100101000100011011011000111000111001011011011010010101010110100011010110010100001"),
("10100111100111000011000001001101101011100001010010101110001110010011001000100111001001001110000010100111001010100010100100011001101010101010010100110011111110100011010011010011001100011101001100101010111110010010101001110010001100101111010110110100000100011010100110010110101100111000000100110100010011011011000101100100101100000010001000110001110101110011001011011111001100000010101110011110010110010010001001110001101100101110001110101001111010011010111000110000001010110010101010011110100110000010111000110011"),
("00100111011011000011010111000011101101001111110110100100001101000011001100110101001011001110110010110101001001111011010000010111101100100010000000101101100101011011010100101010001101000001100010101000000011111011010000101111101011011110000010101100011011101011001001100100001011101101001010100001000000110010100011111011001100111111001100110011011111011011000100101000101100100111110100110100111011011011010001110101001100100000110000011011001011000010101101010100101100100011111110110011011101110010110110101011"),
("10101000101110011010100010111010101011110111111100110101010010110011010000000100101011011010010110110100010011010011010001010110001101001101010010101100010000111011001000101001101010111010111110110001111100101011001101111111101100010010010100110001100001100011010000001101001001100010110100110100010000010010010110011100001011010110001110101000111101110011000000111000000011001010000010110101000001111010101001010011001101010010000000110000101101100010101000000100101100010101101110110011010010110010110111111110")
);

 TYPE fixed_point_array IS ARRAY (natural RANGE <>) OF std_logic_vector(15 downto 0);                                  
 constant bias_array : fixed_point_array(0 to 31):=  ("0010100011000100","0010101101111111","0010010011000011","0010110000000110","1001100100001010","0010010101001100","0010010111101101","1001101111101110","0010100100110010","0010010100001111","0001010001010111","0010101000000010","0010010100110000","0010010011111101","0010001001001110","0010100100111111","0010110101010101","0010100110110110","0010010010000111","0010100110100010","0010110101000100","0010001000010111","0010100110011011","0010101011100001","1001101011111001","0010101100110111","0010101100101111","0010011111100000","1000111101001101","1010000001001100","1010000011000111","0010011000011110");
 signal  reg_Layer3out : fixed_point_array(0 to 31);
 signal weighted_sum_array : fixed_point_array(0 to 31);
 
 
 
begin

  gen_neurons1: for i in 0 to 7 generate
    N: Neu_Ron generic map (N => 32) 
    port map(
      clk => clk,
      inputs => layer3_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer3out(i)
    );
  end generate;

  gen_neurons2: for i in 8 to 15 generate
    N: Neu_Ron generic map (N => 32) 
    port map(
      clk => clk,
      inputs => layer3_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer3out(i)
    );
  end generate;
    gen_neurons3: for i in 16 to 23 generate
    N: Neu_Ron generic map (N => 32) 
    port map(
      clk => clk,
      inputs => layer3_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer3out(i)
    );
  end generate;
    gen_neurons4: for i in 24 to 31 generate
    N: Neu_Ron generic map (N => 32) 
    port map(
      clk => clk,
      inputs => layer3_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer3out(i)
    );
  end generate;

 
  
  -- Update output
  process(clk)
  begin
    if rising_edge(clk) then
      Layer3_output <= reg_Layer3out(0)  & reg_Layer3out(1)  & reg_Layer3out(2)  & reg_Layer3out(3)  & reg_Layer3out(4)  & reg_Layer3out(5)  & reg_Layer3out(6)  & reg_Layer3out(7)  & reg_Layer3out(8) & reg_Layer3out(9)& reg_Layer3out(10) & reg_Layer3out(11) & reg_Layer3out(12) & reg_Layer3out(13) 
                       & reg_Layer3out(14) & reg_Layer3out(15) & reg_Layer3out(16) & reg_Layer3out(17) & reg_Layer3out(18) & reg_Layer3out(19) & reg_Layer3out(20) & reg_Layer3out(21) & reg_Layer3out(22) & reg_Layer3out(23) & reg_Layer3out(24) & reg_Layer3out(25) & reg_Layer3out(26) & reg_Layer3out(27) 
                       & reg_Layer3out(28) & reg_Layer3out(29) & reg_Layer3out(30) & reg_Layer3out(31);    
     end if;
  end process;

end architecture structure ;
