library ieee;
use ieee.std_logic_1164.all;

entity layer6 is
port ( 
       clk : in std_logic;
       Layer6_input : in std_logic_vector(511 downto 0);
       Layer6_output : out std_logic_vector(255 downto 0)
       );
end entity;
    
architecture structure of layer6 is 

component Neu_Ron is 
generic( N : integer := 4);
port ( clk : in std_logic; 
       inputs : in std_logic_vector( ((N*16)-1) downto 0);
       weights : in std_logic_vector( ((N*16)-1) downto 0);
       Bias : in std_logic_vector(15 downto 0);
       weighted_sum : out std_logic_vector(15 downto 0);
       neuron_output :out  std_logic_vector(15 downto 0)
      );
end component;

type weight_array is array (0 to 15) of std_logic_vector(511 downto 0);
signal weight : weight_array := (
("00110011111011001011000111111001101010010110100100101101101111110011010101101100101011111010101100110101110000100011010100110000001000110000010100110001110101011010101011111001001101001110110110110101001111111011010010101000001010100000111110110001110011110011010001010011001011100011110100110101111001110010001111110100101010101011111000101101010110111011010010100001001101011101100110101000000101100011011001111110001011100100111100110100100000000011001110010101001011101011110110110001000100001010110101101001"),
("00110100000011110011010001101000001100011011100000100110111110101010111001101110101101010011111110110000010111001010000000001010101011110010011010101110010011110011010100100000101011011011100100110000010010010011000001101111001100101010001000110101101010100011010100001010101011110001101000101110000001001010111111101000101100010000100010101001100100000011000100010111101011000001000100110100101010000011001011011010001100101000011110101110110111010011010000000010001101010111110110110011010011010011010010001101"),
("00110011101010101011010010110111101010100100010110110100111001111010111010011001001100110110000010101010111000100011010100010110001010011000010100110001001110001011010100000111101011011111110100110100111010000010010101010100001101000000100110110010010101011010111110000000001100001011011100110010100101111010011000010000001101000111110000101011110111101011001111011110001100101010101100100101000100110011010000110110001100001000111010110100110010010010111110000110001010000001001010110001111010110011010111000110"),
("10101110001100010010011111001111001001101111111000101101110011100011010100100110001100010101001110110101101001100010111001110011101011001111010100101100000110101011001010000111101101011000000110110101100010001011010000010101101100111011101100110011010100010011010010110011001101011000111010110011110100000011010000100001101011110011111010110001000000001011001100110100001101001101111010110101010100101011010100101111101101000100000100110101100011000011000000011010001011001001101010110100011100011011010110011010"),
("00110101100100011011010111001100101101100010111010110001010111101010110000110001001100111010011100110010000001101011000011001111101100101010110000101011010100111011000001011001001100011000100000101101100010101010111110100111101101001101110100110000000010100010111001000111001101100111101110101111011001010010101110011111101101010110100000110001110000001011010011110010001100011010011000101010100110010011000000110101101101010000101010110011011110111011001100111101001100000010000000100100101111011010111010110010"),
("10110001111001000011010100111001001101001110000110110100110001111010010011111000001011110101011100110100011100100011001111010001001101001010111000110001101010101011010000000010101100000101010100110100110000010011000010101101101011101001111000101011111001111011000000110111001101010001100110110001000001101011010000110000101101000110101100101011101010010011011010011110101101001101111100110010011110000011001100010100101011001001110000110000011010001010011101000000101011110110001000101110010101100011000101000000"),
("00110100011001110011000010101001001101001101110000110101001101101010111010100100001100111100111100110100111111100011010101010101001100111001100000110000110000100011000111111010001001111000101110110001000100101011001010111010101101000000101110110001001111110010011010010011001100101100000110110101101011100011011001101110001101000000000110110110000000000011000101001010101011110100101000110100011101000010000011011111101100111000100010110101101100010011001011011100101100000010011000011100110100011011011011101100"),
("10110100101111011010110110110110101100011111100010110011010011001010010011001010101100111100000110110011001101111011010000101001001100011010001100110101010100100011000010001110001100111001011000110001001100111011000111000100001100010100010000110011111101100010100111111000101101010100101000110001010101001010110111000001001100010100011000110100001111000011000101110101101101011100111100110011111010100011000110110101101011100111101000110010101100001010111111001101001101010001100010110101010100111011001111000100"),
("10110101110000100011000110110110001100011101110100101111100011111011010000100111001101000100100110110011011010111010110100000011001100101000010110101110110010010010010010101000101101011001000100100001011101100011000000000110101011111010111110110100101111011011010010110011001100101110001010110011111010011011001111000111101101011100000100101111000000000011001110000110001100010000000110101100111111000011001100011110001100100011100110110000101110000010110100010011001011000100000010110000010100010010111011110111"),
("10110110000101101011010111010111101001001010101100110000100100010011010010110000101100100000110100011100100011011011000100101000001100000110011000110100111010101011010110001100101101010100101110110100110101000011001010010100101100100110011000110001100111011010110001001000001100101100110000110010110101100011010010101001001100011100000110100001110001010011010010110011101100110010110100110010011010000010101101110000101101001111110000110000010101100010010101000110001011111010111000100101001101010011000010001101"),
("00110101111010000011000110110101001100101001010100110110100001100011010011100010001100100011110000110100000010111011001100010001001100101101110110110101111011110011010000001010101101011110000010011110111101101011010010000001001101010100100100110000111001011011001101100110001011011110111100110101001010010011001000011110001100101011000100101110110100000011010111100001101100001011111000101111001111111011011000010011001100000001011010110101000101010011000100110001101101000001110110101100000011110011010010101111"),
("00110000100110011010000000011110101100101000000000101001111100111010010001100100001010101011100000110010000110111011001110000011101101000111110100110010100111011011010110100001101100000000101010101010000111001011010000111001101011110101010000101100000110101011000110011100001101101001101110101111101001001011000010101101001101000010010110110010011000011010100100000110101100011110010010110100001000100011010011011011101100011110010010101101000100101011001001110000101100011011101000110100000011010011010110011010"),
("00110000111111000010110010110111001010100110000000101001101011000011010100110011001001011110111010100110011011111010100111100111101100100101101010110101111010101011010101010011001011011010111000100011111101110011001001101000101101000001111000110100111010101010111000011100001011111100110100101000111000110011011000111111001100100101111010110011001111101011010010111011001101100000100110110010101010100011001110011101001010010011101110110100011001111011010011110100101010001101111010110000011010110010111110010011"),
("00110011001000001011001101010000101100110001111000110000101011101011000110100001101100111101010110101110111000011011010101111010001100110111101110101111101011111011010000101001001101001000110100101011001111010010110000010001101101000001011100110010110001000011000100011000001010011000000000110101101100000010110110000001001100001101001000110100011100000011010010011011101100010001011010101100001110111011000001000001101100110111101000110100000110110011010000110010100111110000101110110101101101011011010011111110"),
("00110101100010111011001101111110101011110101010110110011001111100010100000110100001100011011011010100110100111010010100000101111101100011100111010010100000011011010011001110000101100000111101000100010110001110010110101110110101100111000110000110101000010100011010111010010101011000111001010110011001111110011001001001101101100101101000010110100001011000011000010001100001011011110010010110100001100110010110011000101101011011101010100101011011011100011010001001010001101011101101110110100101001100011010000001001"),
("00110001100010011010110110010011001101011001101010110011000110000011010010111111101010001111010110100111001101101010111001010110001101000011110110110110000100100010101011101100101011010110101000101101100001001010101001101100001101000011111010110110000101111010110000011100101001101001010000110101010110001011001110011111001100110000111000110001111110100011010001000001101101001110111000110000011100110011001010101001101011100010111000110011111001001011001101010101101100110110100010101001001100101011001010111110")
 );

 TYPE fixed_point_array IS ARRAY (natural RANGE <>) OF std_logic_vector(15 downto 0);                                  
 constant bias_array : fixed_point_array(0 to 15):=  ("0001010011111011","0001110111000101","0010010010100011","0010010000100111","0010001000010001","0000100011111101","0001110010111000","0010010000010000","0010010011011100","0001010001010011","1001000011100111","1001010011110010","0001011010010110","0010001001110110","1010000010110110","1001000100011001"
);

 signal  reg_Layer6out : fixed_point_array(0 to 15);
 signal weighted_sum_array : fixed_point_array(0 to 15);
 
 
 
begin

  gen_neurons: for i in 0 to 15 generate
    N: Neu_Ron generic map (N => 32) 
    port map(
      clk => clk,
      inputs => layer6_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer6out(i)
    );
  end generate;

  -- Update output
  process(clk)
  begin
    if rising_edge(clk) then
      Layer6_output <=   reg_Layer6out(0)  & reg_Layer6out(1)  & reg_Layer6out(2)  & reg_Layer6out(3)  & reg_Layer6out(4)  & reg_Layer6out(5)  & reg_Layer6out(6)  & reg_Layer6out(7)  & reg_Layer6out(8) & reg_Layer6out(9)& reg_Layer6out(10) & reg_Layer6out(11) & reg_Layer6out(12) & reg_Layer6out(13) 
                       & reg_Layer6out(14) & reg_Layer6out(15);   
     end if;
  end process;

end architecture structure ;
