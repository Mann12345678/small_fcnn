library ieee;
use ieee.std_logic_1164.all;

entity layer4 is
port ( 
       clk : in std_logic;
       Layer4_input : in std_logic_vector(511 downto 0);
       Layer4_output : out std_logic_vector(255 downto 0)
       );
end entity;
    
architecture structure of layer4 is 

component Neu_Ron is 
generic( N : integer := 4);
port ( clk : in std_logic; 
       inputs : in std_logic_vector( ((N*16)-1) downto 0);
       weights : in std_logic_vector( ((N*16)-1) downto 0);
       Bias : in std_logic_vector(15 downto 0);
       weighted_sum : out std_logic_vector(15 downto 0);
       neuron_output :out  std_logic_vector(15 downto 0)
      );
end component;

type weight_array is array (0 to 15) of std_logic_vector(511 downto 0);
signal weight : weight_array := (
("00110001111100000010110111100100001001001011010100110001001000110011010010111011001011111000101100110010101000010011010101011111101100110010000000110001010011101011000011000010001100110000010110100011100001011010110101010010101001010000110010110100100000111010111011010100001010100001011000110011101001001011000011101000001010010000000010101111111101000011001111001000001101010111100010110100100110001010111000011111001101010011001110110101011110110011011011001111001010100111111100110100001011001010101010011110"),
("10110100101001001011001110111010001101010101101100110101100011001011001100101111101001100110010000110100110101110010101110110011001011001001000110101111101100100011000101010111001100110010101100101011001000100011010100000010101101010010011110110101100001010011001011100001101100000010011110110000000001111011010000001110001101010011111010101000001111110010011100011111001011100001110000101011011111110011001100001011001101010111001100110001101110000011010101111110001100110001101100110000100100111011001111010100"),
("10101100000100010011000000000110101011111011100000110101000110011010110111000110001010000010001110110101100010110011000001011010101101011010101100110100100101101011010001111100001101001111010000110000111000110010101000000101101101000110011000110100001010100011001000010101101010110000100010110011110010100011010111010001101101010101011100110100001111011010111111010111101001011100011110110100110001010010101111110000101001111100110000110100100101000010011011111111101011110111110100101110101111000011010011110100"),
("10101101010001110010110000001000101100111110001100110100111101011010110110100100001000101000100010001000010110101011010111101111101100011011001110101101100111010011010011111101001010010111110000110011110001110011001101011101101011100001100010110101000100011011010001101110101011011110111110110000101000010011010111011101101101010011000100110011001101000011010110011011001101000101011100110010001011001011001001010100101000001101001110101111010110100011000000011001101100000011111110101100111011011011010011110111"),
("00110101001010100011001110010110001101011011011010110011001011111010110111110100101011001011000110110100111010000011000111011000101100000011010100110010010001011010111111101101101011011110100110101100010101110011010111011101101011010010100100101110101001010011010011011011001000100011000010101000011001111011001000001111101011111111111100010001110101110011000101101101101001000001010010101100010100111011010011111100100111111010000010110010001011001011000110111101001100101101001000101110110001001011000011011000"),
("10110101010000101011001000001110101101010011000000101111100000100011000101010101001101001000000000101100111111101011001011011010101011001010000110110100101111010011001001111110101101000010111010110011000000101011001001101010101100010011010100110010000000100010011100101110001101011110111110110100100011001011001010000001001101001101000110110101011110111011001001101010001101000100101110110101001100100011001001010111100111010001101010110010100010101010101001000100001101000011100100100111110010100001100111100011"),
("10101000110111011011010010010000101101001101010000101101100111011010011101110110001011110010011000110001000100010010010100010100101101010010001100110100110000001011001101110001001101010111010110110000100111000011011001100000101101010000000100110100011010011011001011011101001101010110100010110100110001110010000101111011101101010101110010110010001100000010111111100100101100110010000010110100110100111011000111011001001000101011101010101110011001101001110010010010101101011001111010110000111000111011000011011001"),
("00110110010111100011001101011110101011011001100100110100001000101011000101010010101100111110001000110100100001001011000110110110101011111110001100110100001101001010111110010010101100011100111100110101010110001011001110111110101100000100110100100111000000000011000101011111001101000110100010110011011111111011000010011010001101010101000100101111010000100011010010001001001101000110101100101110100001011010111010101000101011001010010110011110111011100011000110000101001010101110010100110101011010011011001010111110"),
("00101100101110111011011000011100101011000011000000110001111110010011000101101100101001001001111110101110010010000011001101111100001100110000101100110101111001100011000001100000101100110010101100101000000111100011010101110111001101000000100100110000110011110010011111000110101100000001010010110100100100001011000000101111001101001101111010110100001100101011011001111001001101101101011000101111101111100010100110110110101101000000001100110100110110110011001010001000101100011011001010100011100110111011010111000111"),
("00110100100000010010001000010001001100111101111010110010011010000011000110010101001101000001001000110100010110010011001010000111101100010100111110110100000101011011001111011001101011110000010100110101010000100010110001101111101000101111110100101111001010010011001001110100101010111101000010101110010001001011000110011011101100000110011000110001100100111011000001100101001011011110110100101101001111100011010100010011001101010100010010110001100011010010100000101101101000101001011010101010111101011010110110001001"),
("00110010000101110011010011110101001100110101000110110010011111001011001000100100101101011110001110110101000101010011010001100111001100100101000000110000100000110010110111001011101101100000010100110000000110101010110101111101001011011100001000110001000011010011001110000101101011101111010010110110000101110011001110101101101100100111111010110100100010100011000100111111101100101010001000110001010100011011000110100100101100001111110010110000100101000010110110001101001101000001010100110000000010111010100011110111"),
("00110101000110110011010110011011101011110111010000110101101111001011010000000101001000011010110110110001011101101011000110001101001010000101010110110100101011110011010101101010101011100111101100110000010101100011010001011111001100101010010000110101100011110011010011010101001101010100111110101110011100111011011011011101001101010100010100110011110001111011000101101010001011111111110100101110001110000010110110010011101010000001110010110100111011101010110001111011101010010100001000110100000011101011010001001011"),
("10110101000000111011010011000011101101000000110110110001110001110011001010110010101101001110001010110101001010111011010011110010001100001000111000101100100000100011010111010101101010110100101000110101100110010011010010010111001011011110011000110011010011011010101010110100001100001001001100110010001010111011000011011010101100011001100100101011010101000010011110101110101100001000101100101010100011010010110110001100101001000100101110110100100010010010101010110100001101000010100100101110011000001011010110111111"),
("10100110110000111010100011101001101010111011100100110101000111101011010100011111001100000000011000101011000101111011000000110011101101000100110000110011000010010010111000100000001100001111000110110011111101110010110110011101101011000101010000110101010001001011010101011001101100111110011100110010000101101011010011010100001101011010000100110100010111111010110010110010001100110110101100110010111110101010111111001110001101001110001100110110101011011011010011001000001101100110011010101101010011101011010000101011"),
("10100101100010110011001010110111001101001011110010110000001110011010101111010111101001111001010010110101011010011011010011111000001101001100001110110000111010101011010001111011001100011001101010011111101011100011010111000000101011100001101100110001010000000010111110110111001101010001110100110110001101000010110110110000101101001110001000101000100011100011010001011000101100111010001010110001101101010010101101010111101101001000100000101011110111111010110010000110101011001100000100110001111000101011001010110000"),
("10110101010010011011010011110110101101000100100010101110000011001011010000111100001011001011010100101110101100111010110000001110001010011111111110100101011111001010101100001000001011010001101010110101110100001011001111101011101011000000000010110001000101100011001001110010101100100110000010110100011100010011010110011100101001100100001000110100000000101010111101000100101010100010111110101001000011100010110100110110001101010110101010101101100101110010100000011111101100011011000110100000001100001011000011011011")

 );

 TYPE fixed_point_array IS ARRAY (natural RANGE <>) OF std_logic_vector(15 downto 0);                                  
 constant bias_array : fixed_point_array(0 to 15):=  ("1001110011010011","0010010010000000","0010010010011100","0010001100011011","0010010111011000","0010001101001110","1010100010111111","0010100101101111","1001001000111110","0010011101001001","0001111110000001","0010100100100001","0010010011011000","0010011100000000","0010011100111110","1001010100001111");
 signal  reg_Layer4out : fixed_point_array(0 to 15);
 signal weighted_sum_array : fixed_point_array(0 to 15);
 
 
 
begin

  gen_neurons1: for i in 0 to 7 generate
    N: Neu_Ron generic map (N => 32) 
    port map(
      clk => clk,
      inputs => layer4_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer4out(i)
    );
  end generate;

  gen_neurons2: for i in 8 to 15 generate
    N: Neu_Ron generic map (N => 32) 
    port map(
      clk => clk,
      inputs => layer4_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer4out(i)
    );
  end generate;
  -- Update output
  process(clk)
  begin
    if rising_edge(clk) then
      Layer4_output <=  reg_Layer4out(0)  & reg_Layer4out(1)  & reg_Layer4out(2)  & reg_Layer4out(3)  & reg_Layer4out(4)  & reg_Layer4out(5)  & reg_Layer4out(6)  & reg_Layer4out(7)  & reg_Layer4out(8) & reg_Layer4out(9)& reg_Layer4out(10) & reg_Layer4out(11) & reg_Layer4out(12) & reg_Layer4out(13) 
                       & reg_Layer4out(14) & reg_Layer4out(15);    
     end if;
  end process;

end architecture structure ;
