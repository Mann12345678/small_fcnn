library ieee;
use ieee.std_logic_1164.all;

entity layer_2 is
port ( 
       clk : in std_logic;
       Layer2_input : in std_logic_vector(255 downto 0);
       Layer2_output : out std_logic_vector(511 downto 0)
       );
end entity;
    
architecture structure of layer_2 is 

component Neu_Ron is 
generic( N : integer := 4);
port ( clk : in std_logic; 
       inputs : in std_logic_vector( ((N*16)-1) downto 0);
       weights : in std_logic_vector( ((N*16)-1) downto 0);
       Bias : in std_logic_vector(15 downto 0);
       weighted_sum : out std_logic_vector(15 downto 0);
       neuron_output :out  std_logic_vector(15 downto 0)
      );
end component;

type weight_array is array (0 to 31) of std_logic_vector(255 downto 0);
signal weight : weight_array := (
("0011011000100000001010110100100100110011100111110011000011010001001101001011110110110011010101110011001100001000001011001010011010110011010011011011000100011110101100111011001000001111000011100010101001111000001011011111010110101001010000101011010101001111"),
("0010111110100001001101000100010110110100000110100010100100101100001101001011101100110101011001010010110100001001001101011000000100110001001000010011001011111001001001010111110110110010111000000010100101000001001011010101111110110010010010000010111000001001"),
("0011010011011111001101001010010110110001010100001011010010000010101101000110100110110001001101001011010100111010101011011000111010110000111100100011011010101110101000110011110100110100010011000011000010011011001101100101111010110101100110111011000111010010"),
("1011001000100100101100110000111100110011010001010011001011110011001101011110110010100100000010110011010010011001001101000100010010011110000110100011011000011101001011000010010110101110110110110011001100001010101100111001011110110100000001000010011011000001"),
("0010110010000010001100101100101100101101011110111010111010110001001100110010001010101111000011000011010101010101001011010101001010110100110011010010011001111110001100001010111100110101100010100011010011000011101100011101111000011001001010011011010110010111"),
("0011000011000110101001110011100100110100100101010011010010101010001100110101111110110000000100111011000001000100001100011111001000100100000110011011001011000100101100101101011100110100000110001011010001110010001101000001000110101011001101011011001111010100"),
("0011000000011010101011011100111000110001111010110011000101100110001100010111001110110010010000110010111111111101101001111000001000110110000011001011000011101011101101011001111110110010110101011010011000000011101101010010111010110101011000101011000001100011"),
("0010011100011000001101011011000110110110010111010011001001101101101100100001110000110010010010110010011010110000101100010001110000110011010010011011000111101010001000010111100110110001011111110011010101011001101100111110100010100001000001000010111010010010"),
("1011001111001100101011010111100010011011011110110010011010011111101010111101111100110011000011100001111111001011001001111001101110110011001110011011000010100010101101010010001110101110001000110010111101110101001101001011110110110001111000001010101001010001"),
("1011010000111001101100011000110010110001101010101011010110001010001100101110110000110011111110000010111101001000101100101100011000100000101111010011010000000111001101001101110110110100100000100011010000001010101011100111000100110100100001100011000110100110"),
("1011010100101101101011000110100010101010000110100010110111111010001101010110100000110100011110111010111110010101001101000000110100110100010110100011001010001100001010100011011100101111100110010011001011001110101101000111010000110000010101001000111101101011"),
("1010111011001010001101010011101100110001000100011011000111101011001010101001101110110001100001110011000100100110001100001110111000110000010110011010111101101100101011000000000100110100111000111011010000000100001100110000001010110010011000010011001100010110"),
("1011010010100001001011111110010110110011001100000011010100010111001100110100010100110001001001111011010010111001001101001101100100100101100111010010111101011011001001100011101000100001011001010011000001000101101100011000010110110011110011001011010001011001"),
("0010001110110111101011100100000110110100100101111011000111111011001011111100010100110101000101101011000110010011101101010111111010110100111111111011001000111101001011010111000110110101011010010011000000110101101001000011110000101011011011000011001010011000"),
("1011010110100010101100000100100110110011010011110010101110110000101100111001101000110000011100011010110001101100001011000001001000110000111110010011010000101111101100001110110000110001111010100000110000100010001100001111010010101100000100111011010001101110"),
("0011010010100011000110000011100000101101110011010011010111010101101101011011000110101001100111100011010101001100101100111001101010110011010111101011001101111010101100011110100110101000011101110011010111000010101100111011010000110100000001000011000001100011"),
("0011010101000110101100101110001100101010111010011010011000111111101100111101011100110011101101011010110100110000001101000101011010110000111010000011010110010111101100110010000010110001001111100011010011011000101011100101111010110000000001110011001110111100"),
("1011010111001011000111010100000100110101001011110011010010111011101011110110000100110000110010101010111010010011001000010110101100100111101010001011010000110110001000011100000000101101100000100011001101100001001101011100011110101000111101011010100101110000"),
("0010110110011110101100001110000010110010101110110010111110010111001101000101101010110101000001000010001011111010101101000110010110101111000100101011001111101001001011010011101110110001100101010011011001011000101100001011111000110100000110100010110110001111"),
("1011000100101110101010101000111010101111110101111010110000010000001011100001010010101000010001011011010111111110001101011110000100100101011001000010101111010001001001000100001100110100111011111011001101100010000110110011101000110101000111010010010011010111"),
("1010101000010101101011101000001110101100000111101011010011000101001100010110101100110100110010001011010101100101101100000110010100011111010101110011001100000101001101000100110000110011101001110011000001001001101011111001011100101100001110011010100000011001"),
("0010101010100110001010000001011010110000010101011011000001100101001001100010010110110011111010001011001010001001101100000100001100110100101101000011010010101100000111001011100110101100010000001011001000010001101100101101111000110100000001010010100010111001"),
("1011001010011000001001000100100010110010100100011010111011001011001100100110110000110100110110111011000000111110001011110100011010101111111011010011010101011010001100100101110100101011010011000011010100011010101011000101110110011110110100001010100101001110"),
("0011011000001011001100101011011000101100001111000011010111010001101100001000111000101101000011000011000100101100101101000011001110110101010001000011001000010111001100011100111000100101100001101010110001000101001101001001100000110100001100000010100111001011"),
("0010111101100001001100110111011010110100011000000011001111101101001101010011000110101110010001001011010001111000001100011100000110100001111100110011010101001100001010101110011110101100100011111011001101101000001100011101011000110000100111011011000010100011"),
("0010010100010110101101001100011100110101000011011011010011111000001101011000101010110011000110100011010100000101001101010101111110101000001011010001000001110011101100001110111110110101000101101011010001111011101100111000011110110000101000000011010111110011"),
("1010011110110111101100101100110110110100010010110010110101000110001101011101101000101100011010110011010110110011101100000100000000110101110010110011010100010010101011110010111100110001001110011001110110110110001100000000000100110101010011111010011110110100"),
("1010110000101010101100010100011100101000001011011010110001001101001010001001101000110100001110010010110110001000101011001110010100101110110100001011010100111011101101000000010010101101100101011011001110110110001100111110110100110100111000111011010001000000"),
("0010100111111110101011011000101010110001011111010010111111111000000100111111111110011100100110100000000101000100101011000001110010101001011100101011010001111000101010101110001110101101100010101001110101100011101100000010100110110101110100111011000000111110"),
("0011000000010001001101010110100110110101000001110011000000110010101100111001001000110100011001110011010110111100001000001001001000110011011111010011001111111101101100010100011010110100001110010011010010010000101011111001000000110011011100000010111011001110"),
("1010001111000101101000111101100110110101001110000011000001110000001101000101011010110000100000010011001011101100001100101100100000101111100011111010110101001111101101011100100010110011001011001011000011011011001100001110101100110010101011111011010000111001"),
("0011010000011111101100011100010100110001101110101011001000000000001001011001010010110100000000001001100100000000001000110101101100110100111010110010110111100101001100001010100010100111101011111010100111101110001100110010110110110000110110000001000100101010")
);

 TYPE fixed_point_array IS ARRAY (natural RANGE <>) OF std_logic_vector(15 downto 0);                                  
 constant bias_array : fixed_point_array(0 to 31):=  ("0010000110100001","0010111010110111","0010110000010111","0010100111100011","0010011010110010","0010110111111101","0010011110011001","0010101000100110","0000110111110101","0010110001101010","1010100010100100","0010101101101000","0001001100100001","0010101001001100","1010010000110000","1001110001101010","1010011011010111","1001110001110011","0010101010100111","0010010000011001","0010101100101111","0000110101010110","0010100100000111","0010110000101000","0010001000000100","1001111100110000","0010101000101011","0010100011111110","1010010010010101","1010000111010011","0010011010011111","0010111001001111");
 signal  reg_Layer2out : fixed_point_array(0 to 31);
 signal weighted_sum_array : fixed_point_array(0 to 31);
 
 
 
begin

  gen_neurons: for i in 0 to 31 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer2_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer2out(i)
    );
  end generate;
  
    gen_neurons1: for i in 0 to 7 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer2_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer2out(i)
    );
  end generate;
  
    gen_neurons2: for i in 8 to 15 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer2_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer2out(i)
    );
  end generate;
  
    gen_neurons3: for i in 16 to 23 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer2_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer2out(i)
    );
  end generate;
  
      gen_neurons4: for i in 24 to 31 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer2_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer2out(i)
    );
  end generate;

  -- Update output
  process(clk)
  begin
    if rising_edge(clk) then
      Layer2_output <= reg_Layer2out(0)  & reg_Layer2out(1)  & reg_Layer2out(2)  & reg_Layer2out(3)  & reg_Layer2out(4)  & reg_Layer2out(5)  & reg_Layer2out(6)  & reg_Layer2out(7)  & reg_Layer2out(8) & reg_Layer2out(9)& reg_Layer2out(10) & reg_Layer2out(11) & reg_Layer2out(12) & reg_Layer2out(13) 
                       & reg_Layer2out(14) & reg_Layer2out(15) & reg_Layer2out(16) & reg_Layer2out(17) & reg_Layer2out(18) & reg_Layer2out(19) & reg_Layer2out(20) & reg_Layer2out(21) & reg_Layer2out(22) & reg_Layer2out(23) & reg_Layer2out(24) & reg_Layer2out(25) & reg_Layer2out(26) & reg_Layer2out(27) 
                       & reg_Layer2out(28) & reg_Layer2out(29) & reg_Layer2out(30) & reg_Layer2out(31);    
     end if;
  end process;

end architecture structure ;
