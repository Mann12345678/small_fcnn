library ieee;
use ieee.std_logic_1164.all;

entity layer5 is
port ( 
       clk : in std_logic;
       Layer5_input : in std_logic_vector(255 downto 0);
       Layer5_output : out std_logic_vector(511 downto 0)
       );
end entity;
    
architecture structure of layer5 is 

component Neu_Ron is 
generic( N : integer := 4);
port ( clk : in std_logic; 
       inputs : in std_logic_vector( ((N*16)-1) downto 0);
       weights : in std_logic_vector( ((N*16)-1) downto 0);
       Bias : in std_logic_vector(15 downto 0);
       weighted_sum : out std_logic_vector(15 downto 0);
       neuron_output :out  std_logic_vector(15 downto 0)
      );
end component;

type weight_array is array (0 to 31) of std_logic_vector(255 downto 0);
signal weight : weight_array := (
("0011011000110110101100011111111100110100010110111011001111101100001100000101110010110101011011101011000110111010101101000110110000110010001100101011010010000100001100001100001100110001100101011010111100001110001100000111010110101100001101111011000000001100"),
("0011000001000001101100110101000110100101010111100011010000010100101001100000100000101011001001101010010110101100101101001010000010110000000101011010000111111010101000101010100110100111111011101001101001111101001101100010100010100111110001111010110100001000"),
("0010100111011011000111100001101000110101101100011010000111001100001100001000101100101101000110111011010011100011001101001001001110110011011111101010100111101001101100011011101100110100100010001011010011110000001101001111110000100111111010101011010010101100"),
("1011000000101010001100101110101010101000100101110011011000101010001011100000010100101011111001101011010100100110101100001001001010101001000011001011001110100010101100111010001100100111111001111011000101100010001011111100001110110101000101101011000000110111"),
("0011001001101011001100010101100110110001010001100010110010010110001101010001101010100011011010111011001000011000101101001100000100101101111010110011000001110101101010100010011000101111110100101011001110000011101101010100110110110011010100001011010101110111"),
("1010001000110010001100100011001110110100100101111011010110000000001011000101101000101000010111110010011011110101001101000100101010110010110001000011010010101001001100111000001010110100101110011011000100101000001100001100000010110100000111010001010010011101"),
("0011000000101111101011001010100110110100011001101011000011101001100101001100000110110000101000001011000110101101001100011011111010110000111110011011001001101101001100001101101010101111111010101011001111011110101100000010001100101101000100100011000111110110"),
("1011000000011110101101011000100010101111000110110011001010000001000101010100100000100100101011001011001001110110101011001111100100110000100101011010110110110001101100000111111000110000010000011011010011011011101100111000001110110010010010010010111000110000"),
("1010101110100010001100011000010010110010100100010011011001111000101000001010111000101100001010111011010111100000001010000110010110101111100001111010011111101010001010100111010110110001111010010011001011100011101100110001100000101000111100110011010100100011"),
("1011010000011101101010000111000110110001010011010011000101100011001100101111110000110100100101101010110011011000101101000101100000110010111001000011001001001011101100001011100110110011101101111011000101001000101100000000011100110101000011101011010011100000"),
("1011000101110111001011101001000100110110101001100011001000101101101011000010110100110011001101110010001100111011101100110011101010100101100100010011001010010001101101000111110100110100001110110010110101111010101100000001010100110010010100000011000000000111"),
("1010110010111100001101010101111110110100011000111010111000011010101100011010100100101101000011001010100111110101001101000100110110101100111110111011000010111111001010101010001110110001100010110011001110110001101100010101010110110100011110101010100100001001"),
("0010110111101110001001110011110100110011110101010010101110110111001010010101111010110101000100101011010101010111101100001000100000110010110011010011010011001010001001011010101010100110001011110011001011111111101101011111110100110011010001010010111101001111"),
("1011010101010000001010101011001010110011111010100010110111000111101100100011111010110001010111011011001100010111001001100110010010110001100110100011010011110000101101001110110010110011111111111011010000100110001011110110100000110100111100011011000111110100"),
("0011001111000011101011101001100000110110010010100011000100010011001011110011001000110100010010110011010001100011000111011100111010110010110011000010001000001011101000010100001010101000010110011010110010011100001100100101000010101110011001001011010110001001"),
("1010101110001111001011100110111110110101110010011010010000101010001101010001000010100100101111001011000011010000101011000100111100110001001000011011010001011010001100001100000000110100000001110011001100010100001100000011011100110010101101101010111110100001"),
("0010101000001110001101100101001110110011111001010010101010011101001001010101101100110011001101000011001001111110001011001100101000101101010101110011011010100111001100000000110010101100110111110011010110110111001100011101001100101100111010011010011001101101"),
("1011001000001100101011010000101010100001011111001011010011011000101100010101011100110011101110010011010100100110001000010111100110110110101001100011001101110001101101000000010110110100111101011011000010010100101010001010110000110001111000011011001101011101"),
("0011010011111110101011011111001100110110000000000010101011111000001100010111010100110000101011110010111100100010101100110111100010110011010101001011010000110010001011001010101010101100110111111010101011011010001001100100000100101100000010101011001100111110"),
("0010111100100101101001010000001010110001110111010011001101001000001100001101001100110010001011000011001011101111001100001101110110110011011100010011000110011100001100111110010110110000011100111011010011101000101100010110010010110001011011000010001100101110"),
("1010110011001100001100110011101010110001010010100011011100000101001100011011010100110110001101100010110111010110101010101000110100110100011111111011001010011011001100000001010000110110010101100011000111010101001101000110001110101110010011101011001010000011"),
("0011011001000000001011110101111010100100010000010011011011011100001101011011101100110101111001110011010010101010101011000100100010101010011110101011010001010101001101101000011000110101000100001011000011000010101100001110001000110101011111110010111101000000"),
("0011010011010010001100000001000110110001110101010011010101011011101100010100000000110010010101000010101001010101001100101010100110101011110100111010011000001010101100011001010110101101011011011011000001000100101101000101100110110101010000011010100111110100"),
("0011010011011001001101011000101110101000101011011011001100011110001010011010010000100101011011001011010100110010001011100110101100101011101011100011011001111011001101000111101110110000100110011011010010000010001101010001001100110000001100010011000101111100"),
("0011001101000100101011100000011110110100010101100010101001110110001011100111100010101111010011111011000001110001001101011011011100110010110110001011001000101101101001111101000010100001110111010010110101010000101011011101010010110100010001000011000101011111"),
("0001100010111001101101010100011000110001010111100010010011001010001100001000011100110100010111111011001100110101001011111010000000110000000100110011001101111001101101011101010100110100001010001011010110110101001100001001011000101011100001010010110000111111"),
("1010111110010010001100100100011110101101111110011011001001110101001101000001101000110011010001110011010100001000101011110001110000101100100101110011000010110001101101001011101100110010111110010010111111010001101100101001111100110101001110111011011000001011"),
("0010110001110101101011000010010000110110010001110011010000000111001010100101001010110010111100111011001010010011101001110111000000110001011110010010110011110110101010100100101100100001001101100010111100011100001101001101010000011101110100111010101010101100"),
("1010110100101000001000011011100100110011010011011010110001011010001000111111111100110001110010111011010011101111001101100011111010110100100101000011000101100100101100101001111100110001011001110011010011001111001100111011111110110100100100000011001111001011"),
("0010110100111000101100010101011010100110100110110010101100011101101100111110101010101100011000000011010100101111101101010101010110110101101001010011000101000110000111100011110100101100000100001011011000101111001100000110110100101001011001101011010001000100"),
("0011010011000000101101000000000110110001110001100011010011100101001010000010100110110001110101001011010010110000001011000000100110110011101110010011000001101111001011101001000010110101101101111011000101111011101101001001010010110100001000110011000100001011"),
("0011011101010100001010111010010100101000001111000010011110010001101100101101010110110011010101001011000111100100101100000101110000101011010001100011011100110000101101011011000100110101000010010010000100100010001010111000000100101011000100111011010011111100")
 );

 TYPE fixed_point_array IS ARRAY (natural RANGE <>) OF std_logic_vector(15 downto 0);                                  
 constant bias_array : fixed_point_array(0 to 31):=  ("0010010111011001","0010101011001101","0010101000001010","0010110110100111","0001011101011000","1001011101100110","0000111100101100","0010110011111100","1010100011011000","0010011110111000","0001110010101100","0010010011000110","0010100100111011","0010011000010100","0001111010000100","1010010001010010","0010100010100011","0010100111111010","0010100001011110","0010100101011000","0010101111110111","1010001101101101","1010101000111001","1001100010011011","1000010001010111","0010100011011001","0010100110101110","1010001001101011","1010011101000010","0010010000101101","0010010101001011","1010000111110011");
 signal  reg_Layer5out : fixed_point_array(0 to 31);
 signal weighted_sum_array : fixed_point_array(0 to 31);
 
 
 
begin

  gen_neurons1: for i in 0 to 7 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer5_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer5out(i)
    );
  end generate;
  
    gen_neurons2: for i in 8 to 15 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer5_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer5out(i)
    );
  end generate;


  gen_neurons3: for i in 16 to 23 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer5_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer5out(i)
    );
  end generate;


  gen_neurons4: for i in 24 to 31 generate
    N: Neu_Ron generic map (N => 16) 
    port map(
      clk => clk,
      inputs => layer5_input, 
      weights => weight(i), 
      Bias => bias_array(i), 
      weighted_sum => weighted_sum_array(i), 
      neuron_output => reg_Layer5out(i)
    );
  end generate;


  -- Update output
  process(clk)
  begin
    if rising_edge(clk) then
      Layer5_output <= reg_Layer5out(0)  & reg_Layer5out(1)  & reg_Layer5out(2)  & reg_Layer5out(3)  & reg_Layer5out(4)  & reg_Layer5out(5)  & reg_Layer5out(6)  & reg_Layer5out(7)  & reg_Layer5out(8) & reg_Layer5out(9)& reg_Layer5out(10) & reg_Layer5out(11) & reg_Layer5out(12) & reg_Layer5out(13) 
                       & reg_Layer5out(14) & reg_Layer5out(15) & reg_Layer5out(16) & reg_Layer5out(17) & reg_Layer5out(18) & reg_Layer5out(19) & reg_Layer5out(20) & reg_Layer5out(21) & reg_Layer5out(22) & reg_Layer5out(23) & reg_Layer5out(24) & reg_Layer5out(25) & reg_Layer5out(26) & reg_Layer5out(27) 
                       & reg_Layer5out(28) & reg_Layer5out(29) & reg_Layer5out(30) & reg_Layer5out(31);    
     end if;
  end process;

end architecture structure ;
